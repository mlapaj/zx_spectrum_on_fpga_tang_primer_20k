--
--Written by GowinSynthesis
--Product Version "V1.9.8.11 Education"
--Mon Jul 31 12:55:46 2023

--Source file index table:
--file0 "\/home/cod3r/Data/Gowin/IDE/ipcore/DVI_TX/data/dvi_tx_top.v"
--file1 "\/home/cod3r/Data/Gowin/IDE/ipcore/DVI_TX/data/rgb2dvi.vp"
`protect begin_protected
`protect version="2.2"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.2"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2022-10",key_method="rsa"
`protect key_block
TMsy8SxpC54gwLrtR5NIV4PEq4A9JM52Y+ee6vnooPK2VjnLdVqLrQt+Zcbmp0s0I0xr2f4F8M7c
a9SGm1Ln3bscHZd597sb3czt6bWWTwYUvMIJF+51qREKpXaNacF67DDsI3FaHvOBJNdOTdtk0dj5
9o438prTDR0aRuLUWtr3M0yHQH5PLhM3jUtRH91jiJlYh94bR+wfeva707H0FiExD9AK/FweJafu
La6nOlye6fyju9cMKwLwOyU22Og7QvokjejM7Cq3v2mh/mk3PKHkQ3dFhlrpO/Lc7sJLMcbvuK4c
jOPnd5affrhraeXK7k0NCHOJCxQIi3P5yyv3Qw==

`protect encoding=(enctype="base64", line_length=76, bytes=69408)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cbc"
`protect data_block
wL5WKmcDxdbGXmZir6J3DFgW38vS7n0AdCrsoH8MANJfIzF0Vda5XPI/zG05Y+qgign6Gq8Lwzrg
ncagItHon5FUCZELph/fDXks/Lk32FySmcasimAkPlEkGZ1U0ZnhHDseTKBd36RW80LDJqaHYObx
Lj3wEgci393HUcn+/UfLqx67hbof/bLfyoqJx7lONv8Mqr/bbDT+WaBWUFLj+vb6CzRuuVb/YvZg
K8ijGiphggaGw0Yi6FEVqbydh31UUsDyx16Cl+A4AvN+6W6rcRzSizAO6id53nunXxdtfuUelt9j
4juOgz1zZyS5C+yh1CVFMd53wd9znlseOkoWPhCn/zE1c8VswZnkjCcq7MkD0FALhMjXtF2rR+7b
FDtpIRHLNLVS+d8jAjE7TYTvvIayFnjLytYk06EakQN8rDJGpjt0VORjKnXNEJB9BHVA2bmIgnIg
P6ZR3xtEBdTsUdXF0vqvU9gX/qOGA0dsSkCiYW4fEf5/QQHBiX9KNgPHW2QAMJRBamwjl3357K6O
dCv/Y9ZVFZvQ0uMikNwOj9eGvjeEHKdI79IaNhirOwUoM7/3b1KJFW0ZVkOdEa8ANtwTCiHMXn1P
/OiVoaKwUwTEN15gkV+yxobCNEhVaMA6vcDR2IbOPPX5fN8rY6cC2Lc3TzlxwvYNk5ucFForknMl
OBZkH8TMVWaDTLoSvk6cECDuUNX9aaV7ShBqMHgn/2oTrKD5K6m+ZDJ0avFmMseCDb4XPoLUHxKy
xAPcr9SvQ7SbynpCSzQ8WcWAh5kg76za1QYdhMcPerxOnRzlxEisuJCGDj2DGWNkq1Yr3X3pGtMN
KR3QE/i6pHqg0vftCnn9tFZivQ9vkPCwmJJ4p4T8adCGU2Ru+1JHHUZzxaIx1An2LLFgSyzbturc
99yUu9HcLLxp2ZDhD9QAQ/umsXMhExOXO8iyRgqQvNqmI4Zts8MIwwBRKL5NxrN6u3suxz0fscK4
8RJZgsshCUeZZPn5Y4N3LXM5ysmZkd7Y6LFipdwv5M+ZdCLAb5buLQPWVZHzUKiLvMPYqekBeCRD
5uFipLD32atNzooHhguVwqYockBtZ7DTAiizMGfvYgsFVas8Y+Sb1n4uEMD+QX20gVjMW4l8KpwR
YEi7mufk+CgNMd/3HJpwnISuvn/gOWYPLXNXJeTOH9mqMfqZw9kGCUIPRbzk1zucBobe/sP9TXen
3AAUS0iKU69mNJDiXQDyGhB46FX6vmi0b2yqXzfOUrPFxREFcEd1zBH0eefShIA7Wavg8gayt7Ya
a6E2U7Em6ZFM+AeOeUh2b1ZQAADLTS/XF+tQ/70+5EOBhvkuoUOw58T5vO3KcWCQnzJCeqkCNlPZ
BRWrc2qB49zQddgoWpOAZE1QG8dn0kNWCxp82Btcad4JyBFvRUTwugEMWyGBfX+lfBWutu7ny8Yq
FEI57OdfIokvvmiHCutsNiB+TEzlAfMpiiyYkRZ7c1k5JFPt2IwdIPWmgpPqSFEThW9Cmpqcl1aU
mQGmN1tEWKeKYIjzIW9CxnIK1SA2R1a3zquTobZXzCEH5OdUQ8EqWCrH8usuJ8Y9S+XZYNQ2rZgu
vVy1uhN/oDPWrwTcU5hXoseWVpZHypjrBDJZrs03BbHh9PlZjCpxS8nMY2N78TOoRLuVt8XWP5+P
WEKApjFRPiZvGcWMPXF0nnAb1PjQjWNeyGfiZK8oM7r/rejOJLfcNINO6HY6GbffeCOXd7zZwss9
AZTEjSz2xpKOR2QLrR5Sl8mthlmTseW9ihFUbrfw24+zAU4Jv8MTrgjZTYS53H7waTmK4wN/2hUj
vcLgj1foMf5sgII1xjEDkTtrljbXHfSE9KiC4wKVZQGMCN2WaBuLGUCx3Me6Pe7dgl5W5OZBP57m
7nubEW8CBbbDZtcfiSOUBE4P9S/l9RpC9NHtSYUCYT8bKcrnC5qpE0+HIrpZVDFD6STcOfRbI1k3
ITVPwbFEIEmqJP0gZxlHYxla7qefYoooECZO6S1rW7N/O86NAF4IvhLb+7xA4OR2WrDd7MKjw8gV
o29yfGIbrnRDD/5VIo68fb4MaZNEDDODydQdFLYS4rFKKOa0pmBP7sDYXPEVs/HsG/P/gzBkqx3j
EqQ+4j1RSkHD+besrdmlAyXV6Gk/Jjj88M6A5QntQYxTATmXG8/bdbERNZc61M04DQRAKpBJpacl
WEuFP0pbpu9alFJ+OdPIreq18mhzBt8o5zBh94BfBWg7R5meR+6sB4pLDOR/chidpJgH3vp3GVgR
VmStkM0PZfJheiL5Hoi+K8gEzrFnShXr9q09ViTKJGs26oSTMUvH6XdF4lA4S72jIdtZgFWR/LwZ
UF3rxsO8eCL87rqmmVG3nM84mOYDKtwa+0cJZX1lHWh+h04MXkizQkfeiNQVM8NFC91EEaJCWjQ7
OJq4fzeDlpGLiqR4BKDAEnL50ud+35fJzz0cJj06jP9Jy2T5H1gdsyUVZVSK15bu0ueBA99MVdYb
d0MIQ8HO1QHwlvor5IY/mdPqze1QkPTyZx2vgYqC7GmiHAmh0oOKpfdb3uh6xC5iCQZvZFXx0+3R
D2fCsbmNXfJwoXhJKviZc+tpqPELpFoCql5uTWbHyeDJunGRNs2WvICPEAVXEr4bYsb+Mv2anQuY
EFhtpCmkjYAqSDGS2MUMIWsw9cVp25Ei711y8tt/4nPrUgoZyLEdnhH2ogl3wKOFcs4/NbQVuii2
z/nDTN3OtgLJ/PPR8MBpKGquPtaNb4JoQp1mJvdyBCmggW8cjgkZy0uk7Upu7M67b9no0dI/1uun
FFYlRsc6uIajVzVr7aa+Ark8o470c1txlb/w3j9ntgXr2HBMmJiPXL6LPRF/mpaFQnhxYq36RSwr
b1kkhPhxnpAYL/eQKqiEFkUwMa2bz4/jhhZ1OVNSDSG2eHbHpYaUPQgG/wxx1s3dNmYmrN/sPoJr
LW9SKad5wbOZrbzMXJZHlsWIjXigSTAMtpBC0UI9X6IVvJ3eeZu4moFlTahy6Ak4nNNYAlGPdQgG
kmJEUWQZVe6UNtZHxpMJt+/9V63W2kef9NxP92Dn1w1WLdettSPaRwF+W3TkqPV4LLcuQp7RgDXf
hDj7+87aIBDkMayWcU+V05UJYvfStEsOiKLNTQ0TvdvD7s4Cu37KLXVukAuwEyyQ96q+aKHk5lLA
aeAKuVlnGv3sdU0zJgrxxgz6vljbyCadDauLA+7ZswDMvRWMroJDEh5yOQOTS5iztp0Q5Ca6thhh
uQEz4rPvMA2hlYZ2MzayGcK0DNx3BEkV3HQO9S6lvbcs55IrIR8P5F0yWwUMXYPCtYTZUTvD81Fd
p3YFhEEXhe368uDCMrDApUUFTXOz4weiPzbdRfeDTsajwdZiSkEk2q/hOj1HU0Oh32HkBUKxhDHd
usXA4h9iHgdSx18iT6mhVzAZpLUK5Cul5HdgPuOKLzi78dV9vUrsL5CMYjq7SEpIDaLRYaEbh6Yl
t61tAxfZpbaOUzWenHmAO77xbLxnkTvXyc3r/goikAVfbR85SoUvvQOYpoUhpbv2N2SGjydrYnX8
+WPWKFjJMf8f/q41cDOcy9OnhWKpLikMs1iE+/IcjF3CwCS6LV9K1WEUagsqG4DZrZyGC+S1IoXm
lQFe7ehV9eiC3TnRPgrRhmTZ5cQJAX2tciV0w1b0YOvgHYM17AjAiIFRXHI1pLKhyVoCxiu/f70H
bAQmI6RASZeRzt/WCx6NvQ3CZ5/ghRfcJ1N1Uh4wwSTG11UG+pvT5bV2v1PsCdJB8psJjNYv23C8
HUEk+N8yjkiPM2y2VbA8+1PpHk/o+R20a6QX4EQrnahlzQWka6iLxr0O7UMPi+UsFYEwRIJ0aCcJ
cMspbaNoMReimgqKVa0GFQLm2aqy+HOu27jMV2wb4trPXiAf3EqLQXE0F3iNiQdV68Pe4YMI3OuD
rV07GNa5F1gqmYPjq6D5dRQgmiYqFE3h+H4TuO8jJwji7PjbmLHXWNB3IDUrQGxK50YECAx4HEne
yHbzcqJx3PoYeAIzpbvNjM4ylwBuqFJxjcS+yDwBX6SvZpi85CJv01yrxb0TBIII+41v/ty/FdAx
o1OMayyPhYsjBBbScxePWUl/36u3eqh5JcPTK1Cx8mBqKTwzXrm8Xe+Tchfn6hR/pODHsSlXEQ7z
Jl4j1D8YQFhw7nv+83M+EqJZ0+Uscf/Ac7Kn0ci/PIUb9axBM8HeLppwmtQETtcO6Z3fWpPD6sAy
SWJbDx0twyJdTnB7mbOeQszsfbPzy1FDZG7NX9xb8Ro98LIQrm4BzVbgyOYQHHTzufEeu0nLYdmC
mW7l5Wrtr9jPIp89St/F0aXipO2J7eqDxefKRsqRN5yg43tFcnWJMfsDtDGxTaTLeZQM4zkIjDBK
AqgIMQuKhB5q4wzgPgCJh0NHjfNDU5WmnFQmaf7xyHdn9Hm4jiCStqtlTGx5yGwy5KhxX9TkutXc
PcEguvGT2O/hA4Pu+ckR5KODvdRD4jqNvS+MPE0l7ud6bTp04wsc10DyraMWNs65ofdjlnAi8NOW
rFGO4Si80fKWLU1T91zihJMLkPK0upud/8lfnONpvf7ql9Ar9s0flbYa4q1OIMRH0z9HovdTGrlf
0zD5Io1Vly07awACPgIBLWhyB/w26vIWJI1jQw526PzK8s28XnFLfw345WfCeJY8pUwCHCxWOO0y
sQ74NAzXc7L+sMKU9pcVhQVBg4t4xMd6r43Osz4q9nRUcFY03PApmr3k3tEZv1weqFl9huf9IugW
9Ye1Qa+oOnqaBppf33NfmUn6gLt5uJvDppQ5tE1Argjmvor/1n2Tcp9m1UX9hOL88GqfEfQlc7FO
b2MciGGWD32C1vHp4Bzj6ttoOeRrlm+DxH1HDzz24qV+V9aU3YnaJW+U4s/cooyNFqQxtX4UNiUl
CltlMtSj/TfhprY2Al6DeDxL8czPUdDdbrlPTzXaO+Le5260Xfj6PpxYQsR7r+YOQGdVq2i8MNTz
67iP3OnNcWXgh2zGZclmL1Zq56C/w++/uaW+lhuApp07zn4r4XgjHGqLu7YvFT+Tpllfl4+Cym0+
eHmK8eXmZ6h43/X/y6/o+wdhtsBZxDrLqaLU8US6R/2KuBbaGBQuV0eY3esZ+LsB+cDGpQsb7NSO
Bjr7IhCoZuszb22llWOeZmp0eGXn/5EaFCdBLtP+PaRQSo6oWdNsSMQzu0NclVfO/htUFp5XF3g4
cS1SNOhBVc2VQNRWtR7hJHiZQ+ZJCUNLr5tAzRaeUQ60KfKr7aij+iutUxNnkEEaz9pj81wJMgkZ
mAcQt2Whr+UbJSs7kA5cp6dTXunYSiugMvqGlCbCZvu1yAuosvqYE9pJhnMVuxhQ9BS4vu1bIKlF
JnYadclWKNci3d57DwJ9uV8YwoDsqZ8bZHRKkbYunQRcoP2VrT5ysfmVD8Dv8oessPCINMX0xiwj
FysZHKc8EqyWgHy4YrY/JxLzyzSMTcAZikWORA46ImSeolrNi8OIqV+FTSuhdp6dXjV/ZjoBrihM
dpkS7+RaupEYpKyT/ZU7l01ERaQpmX13KwTeYm6rc5DJRRoMs3d9U5ve05HQ80O2Z2mQ24kf3NXl
35lHDc0sBC6EX3uPI7KiMD3f1kFSCZhW1V2uoQ3vClNZl+Jn0pFrsCVEgPjORCsV+JyPatqZ6Dnn
RGIybNFvCCwX7MFVUs3DA3qOY2wp9me0YdVE5auMS9hrioEp/wVmdpT30SlGU4JL5BNpqSBuFjGH
l+GIWmR0eC5E8rAxGGqvTTY8AirjgLCg45cCbE+ZZ40L8YENrIhzPWCjZ7t9zFM6H4ituZ03REuH
9roR9/i7+AC2qSysSpp5evNn6aJags58GBRJF36g7V4WTvCr0NMj8YhGidLJafxmexE6tQaP85dg
m0nh7ciH4NGy5ebaRsG7z/6xkMn6P3JJpISp8WAWziIni4w3Q99qsW9CjAEP/QxJ6TlneubqDjIw
inzufSOmvMAAWf4u9P+JN39mMu6/CEqERsbEP1/ku7uswjVAJWWmxRfzEM3Aua1sLR9BpiSpkkdL
yYA6/4BR5JRfMRoUph8gpOUrOjSID/lgTwWF4d+1x0IQ4M7bOi/XsuOEOjGw5+j3I98JsUj6c5za
wsyyNyIYCTvrok5oEUk1duvxK7opSVZLfiIZfU1tqjsYeIrUINoF65j0Ik6WhY1MyBwt+jKwsWX9
A/OLJqm+8wFhOvdPTazTW4RtGKZ7pbbxD8/eqkZDynGDXN/cAwc/+4idHyOMWte2ntPfrdsxphtb
HW03BKSU6GuzQrDXM3658MhOI4aGFOppBeuy54hnnYLAU9qy2naXkwlNIU3/yq43qpXO8xXEbNvN
oPTDUSFphMkm5RtNGOgjwBmiIt0Axk30BvCFtNw0zX+StEohojMdcGCd9UXeOyvNXO6FZ587XKSC
wU8f0H3IBfFOPMRkaN9sVbZ7W2Rjwhy+F1o4k6Sauwi+DZfr467IxAUgCheriOTWu1O2OfO3vQ7x
uf6icpG1KsJpVG82D0YxJ7jbKhIf3CEu7ig0yDyWrqvs15gkc/2cLl5AHz0mUCwRKgDmRohJimvO
h8dxOettYwrXPQiIVxxQ+upBik+wJYO6/P4/S8fZ2yaXbjpwBzC/mQminApmn+J8/v5FjVSiLeym
fPyc/Wqv/Sk3Ayj3knj3NayY1alTPxa5BbRns9JBfzy7AyvBBd6DX+128Clh5l6HpZG+Heyty6VK
YHZL0Ccmroj8Ogk7EMC0TTeo782N2Eqp4G0bruGykDe9SVB6bxDxisoSOpECld8MCscHyqYdZSpe
Eq81iNsJnodT89YRY1LmJlkjixKElcVZrgfz8EWscCqY32egnvO3/tEd21XPPN3e3W01S1/n/D/0
SAT7hYBf14baf4o4orv8gwMA4jCGJQCMt8cK9Dw6CORLd8SyAimW897AX6XxcWwtQgLzJSZ9OWGN
/SzHGmHDziwgMWzRCO0N2tmc3Ay07d3pdoiq5fpceDh88HDOVICI9ew+Dhu6ZqLTNbBtuL4IcBv2
QP6Pn8TKre3KMsZINXVB/ui+DH/OC3wnmdVLGK2S+0pbqrKJspcnQ6V9ynfEvqNYm6hHLV9h5N0Q
grXV6OQ1/eC+9OVXOOezGlzEWAne07LKqXaAs2+gwZ03NZrLYFV0oZldJUL/zu7MJrs/ex5KBdaZ
CFhXxLZSEyrnCXlFuDkFibVik7rHYghAxxpnLdKwx0K43jhcn69Lr7O61wLTO1YDzQHJa9TzDDUX
76veR+b4je/QrIM2iZOaTfHGh1floa3RXNUtBPusd/t4CXTNlig6nU99/Z95Wgh5miflMhfcXI5r
is83q3OQzVmCnKbM06wV1uuVlTBGvNAYIcsSGWLmG+7wbQlQDbchvlGRG+ZOaWvQBxBCtqddtFVe
f/XOaZgWeBvKlmMLxfJGAm0o7D4JIpwtVkKtZFj6jeblwCS+1iSWzRcFcp9lSmc/xEWexruCOBTT
T9f7qfhjFifi8Q4/QcnYAgaFD48DXNvINx79s34mRsrr/SsuBAXW5PlqbV05PsznM56skk4M6Ilj
ibd4evhkmO9ZJgMEiGfzJMxTqDk7naj4C5BMOovUwCpIamTsBFffpBNoDr6eMIxTS8oX8g1hvzyH
NgJkxJqfia88Ua24G4n1gicdtfDsbFIYDP98Us0QkkD9J9kbDozsqij81L9VnZvXcctmAqNEt1p5
4pD5SL0+fuoxtbB+QSQonIHCKD5ouRyzmKY7TLdzwUi7nKAjh+usZocL4oWMGkuTCF7WzcgN0yoR
JoHrWxz8YE2pQU/Ke6qYXD1g+IQlGWd+BgQRL8f//IpzzYI4F8/XwZh7bPW6EHZcDcheh8AiBz+2
8OS6x4XPVPjT5rQgOTjzxbtzK14x9DFL/vOF62iFFdRSha2239ZmrcwhHdAaTG2SY1HIkk6ua+/L
o4dhR2kpMMpH4TqxHVA3kksfbHfV3y1A5U/gmpSNzxRFAi+8mYr/oDlOO5nX0T/5Rpddd8q0SxFK
LCe0EJekDplKORGoRJ06mLK40WUdEMOqI+5ATi4cZN3GxmWJFZxxfFBEeS8TOAE5qCE9pL92LNhm
Z2GPxOx/uVAMKrK+esK9krwVgSLnBgpPcOG84PYFlaYETB+FpYOCeKETWnguOVWwYs9iA6dQfbwb
Qu7IlskdXTCq9LEWMGAKwUioUneMHgPLZpDnE7IVTTOHfjAa6T0Hz/sSJwmY+MZt+K0eozIXyJ2F
+yHt2ZbmR/fOFEoRm7VCnthNEDzs4Up1XerwqxkTits+Wv1OIJmxWTIwZEbNnIwJdWx96bQmhXWX
gjphtItgGe2Y6U7vc82vIVMDLtSR1sKnX4ifLcwsveHScMunnyEoj8TICIUOjfkdGypc93jNqzU9
BIEept2Z/3/3Rffpqt4fPb2RPs4yPf6HQZTCzu18AAGu6e73A5igRr/FaILSCE6w4drJt9cQeuFK
syFHoql5nPrcEmqDYJvs9sqL7k6Wg1fBU2JFZ1jSI5nGPn421pYElU3+bptdLt8894FaMU9qKtRe
nHXN1dc5694c+BUygKYzkL/bOvKcuUt96bKGrUiHN5ZgSi096fzrzXi03bPIgtdcRKW04YUQoJHl
wQWl65O/4iJiDfXPFygLd870k8dObqSeUsZy0o6Nti6pBRviTv20wpnpdxJRLzSd63iEzEWQpE5L
C0jI7gXbjx9TFnKoVWl7WlrDJgTpd8Kq/ku8hmwXfyg+NhnxhZPHJqLu9zHiffU5KI93RjGb10VH
KPXb7Ye4K3GRfkkr+Uv2bjH0WfvTlSuor+LAuSgpg/EpCWV4VSLR5tW+kqGNZiacjLXaOJGkGoUE
g6w+ZAM6UeEs8mgsuIWXN2Dza47avmfqoJ+RLC3v5h6UIwNClPhz7SFVI6IT5JlAXXiNcBmqYXNV
BBVcud9a01CjYIms8eWw9iagFZyRGBOUvsESeB9qSzc1UxmZlrlpBacaLMDQSeZ1BpXZZyTeqDvx
B4Qua1kjouHWYPfGFzbjKy2xQq4yxDRqFZ+vyWJ1qIXrahmGxIKK+tMVnWsB6MQvrwbSKT8/n03w
hD6DvM+g0lvfG0tuQ9eThLu8S2LeYyzC4DcPG8eIyT4SPEiQJyooamqu8RJFcz1SkMGTyCHBJKrj
FQp20CIaGCVwGP5R+zj3SM7SXprFBSNLiuossuP+XIK9MI1f+/mXRGFsc9ESJ0uzOZj13NLCc3Br
IP1mriGQfBkDlTIQA68CVmg7V63Q4wVQvNF3xx0vA2Yf9zdgDckDZFqNEVft1eJXJInEs689uk17
cWfi72pu5qQ9jLMxGgtPLhGCPAR/+sFE8mnbw6lZ/rgh7xD4ysQNQzQCsxbwKwaabXkZyitGKIbH
FQischH2bU3gXRn+Qho0ETxZ2SJKCbgm7ZzR8gSR+/kEoRebxzqSet4N8mjy85HmxyaGIyqywPj1
hl8bk9SqXf0TXCLEo3Nr5q19VPk/eYF7ld/vACv1ceVq5pmn80SMnjEKbzqcQCeuKEGQN3/KC/uX
mWjz21R/J/6b8G8TaTy2c8tvz2XukGxlRB4TdAjYdKdEhU5WBs4B94Cy2sMs44otRYsxTpgg1pVy
ffplhlkWxnaSTSNijymk3LqA2gWz2dVm1oWgc5UP96hYnBKrdTcs5YIKx2ibma3MSRellS+LTAI7
5irG2iGEpzAj9j8Xycz2kRrCqR1Bsiz79ZFJzZ2zxP8cItP862IROHISmh6YeFehCi0Jmp2of3m/
g0rop0g06Cqvx4aVa6dXnnuBE/U9EQTXN3+AHGbIk07Q7G1lJsBXRnqPVmmQFoW68A0rAnq6fNUw
CHUYP/EXPyK2kfc2853Ebbjf0miKQ8zxkqZRvFmGR3j8y4Jshh+m62h818ts/ZMCC8Lh2ClfchD3
ROmabBsWkglecq3mGaQ39S/6dKzEqsbWCBgPqW2f/63YhM355j5iyB35NTBTpxR01kTDMtkEA5UY
mq6cZG2lKVdM9+aJR7HedQUGLCS+EjVZxqR5uxAQZbiDHAiyJGoxMsI4j9YtM426ZEgdgF4j/cXc
8XJ/PWpl0fhFFPwGw+OUX0npAOz0hZxmJSpdpbRS+ifEo1gLQJnVpeTLlRpq11fOuJuDiObYpjxK
IyWnu+5ZJ9lqjk+T0obMD1YUySttbnlc2jhI5NcYGtG2UDTOEFaoiw9NypJBcLc+kNn8J5m8JbKP
Q0QioSpO6Sy3Fo1B1NynlgeLQRLBEG8Z1KXJboz99tUcKfIPkt142J4DDFfRWw7u58DN5CrUTR7l
TaY2ZwLiTxn2AwGHX9PdU5EzNYn2kMhc5dUOxZ+TYc8Y6StK8Rj/qKnTSi5yhLNWB9kKVUr5jd+/
qCrgkZ69ybAYvf7pmlBhRMA5vPWgBlr//CGM/AIkTW7HSU9MKjDiUKfGrkOQoPKkgYSyVMpHgZJi
nAoMaKUs7WNcJVgrrMLlGwCcqAYMc/3TP0R5/+fXltdg5gS9noPIUHKTSL2h2RX6VqxvvDOnnlJe
bAVkYc3z8lmMHEnfd2zCYLyp8aVuTriNQKbmkPfl89CxTgia2dstZ99Op8/zGvhtoorRvY0/BZjr
JIaQ3upBDZWuP1f/BWUTaG83bdcHD2Pva6GwTaDhpenNfr+Dp/Hxxe5xHXGdtX7sjURASFW9W4xy
SHaYtWOH/RVnwgkoJNNKqSgBqn+q8lrcBsRfCUC1BdfMhk3HP0vfVx/syDMTyi2V6gaoCSWRpaYh
yPM32qMYtqKe1a26JWp/J6+C6pCN2yjzreKqW/WzL7/9TaFlNhS9gKX4KDSk4i2l7d+AplqV2vKb
7TS+MYIyy8DE7nbZ3kfYjre2Qio7khydliDmpJ7Ds9ibJIKFElefNcRb/mIxV1c7KegAZfLsptxJ
3ZdAHMoiyY5esNCJbHp5EIBcQwRidV8murCtvxGnuWDfPx46BSNC7FJsgH8ezB2XH9YgRwhDrgyn
uvR8qzijbXHVgo/xGEfiC6rjUwumvM6MnV4B64rAcnyWfgpXR1TZD+B+7kkXBSTjQti7h3SUptab
ef+rGED/SkjiDp7Z2NMBhW+zyN2owqK9IWIfkWfD1m0zfPggkDz/XKOZmFAJLVeHxNCj9HQoDubt
mrqAxJvHpAr35SE21K6OHmQAS+zNc34kPcgx/2b6A/faoOeKWGY44GgrYAEII595BqgD0jXXSQRq
X559c9pq5fNF6BLtpiid8vDl3MqWVgUbzb8ZwKucGySonSD8+3ZwkeiItnHnGiFu9lkZrU7mu9a+
vlE/da3f9HKU4axh6W7azqVP1QsceMNZGKunABkB0E11jNI7MA+VrIxDzhJgJDH6DzZDXN4Z/q7q
l1xuRzcr7cUVycWsPBpVCWVS59xBoZHcuuPuQfwCgPzjmHNbLn2nTyeTZqQ601iGwbe10YnJtdfj
FwhJaTQ6gDJRTj980BEIB16BIp6Vs1wTQHMsZeZaY+ZDCAWMzTr8HAxJboFrbXTvT8eKrfu8TEui
gQgrM+TV7rzp1Fk/tTGDf9ClvlGuyg51lKI5MqncfUPCHq7qedG6CLgvefmgv33oWhCUswN+xdKZ
PWRPpbsjpAGbnITXucTpqP6Uuh0nicHOtS9CkZH6tQOWxAgadoiVxpYhWcegX3f1y/fjZB5HCVQ5
FcqQkNpH+OLgQ3y6YudWITV708LNg5qnFkJxmApidfVHYRkKtfP0xpZpTKr9C9U6Q6vCimtBhxok
zdHmN4DXliKUHFtkLaSNQeJwXHgLJszY6rsmAy3x2NAQY7OlVzIoegl5+u6aAvuNR622JSNdIIJz
0eroBoAnh2mgRkqYVmfuQpaPbnjYpCXDdr3iuiWovH40aR7yh3WVdjUjbNsJ/CldyVFyTKEsi4Q8
wNhCIfWMrKNGxvr9ktuivz3+Ym+MqXzZlEUGfBZx1ygGLqlDXtzbAMZOn9F+xzZFSXhAp4z4FlUt
Jfo56VfiKGTwKN5I+66zTKp9wibLFZnD5u0RKkTm94dJEPoY6NVXorcQafWI9isfy51baZ9VNrRB
FrstpZuyyv+Roq6Rdm5NfUCWFbklrCnUwytZUYzni5WdBAlLOHBJzURIGZVIy3YwS1NGzX/MRz8z
tADbUux9U0VxtL8eWIOTy1ML3o24EsH9ZsqZj+zqjsfm7CuysbByo3jdQxLiiHlJANF0dnrVy0nb
5KH3EteZZM5+BS/c6ydoAi518C6iUr2CAQbL6AjDMIAMZ/RyMeih189XuHXu3I8aHCRSV2f0VFte
4ILDyOxplvrKSHJSHK0a12SiTKuEVKJXPi/IXlzvGSUWt4vX1MZxAgTCvlyKrXo/6x2C6HIUEQ2H
olSgAkIjDaiYcEGy7hgZVxIcUhJk8eTau4BW1RpoSsGYwOGa2XiD1RBzwBcAwR04CUV9VArhHugh
y+O1mldDR7JkE1GD+88y7Ui3QmJgOfs8Hz6gt6fPLqHEajJc3Gf0pZFk5OcUjUt3huvOjuvBRMFl
ZbhvwvGpuu2Hkx7JsnCnPJkxHJQXOG81Hue70tAye2wCmPygVqfF2KYxwZHu92EidABsUSNAkgMj
PJAW6U/+ks+yIG2khu4cA6Y3vPz816/VP8HXeyR4D9zQL3H0TZGdqSHTkSoQt4AtuHUwm04JkRZN
cddq1zgK99as1ma2LWxAUaBKCEqF/l1H1V283HNG0QRZnIeTjzaOIJwFJDBOHHAqb9v4YrdpviOm
GbEvPr2UvuWWW0nC2mAFqYZxbgHMkcAIsBxeaRPHj/VP1P7hLiV5+wUFaDStmCrb8cEgPLmuHUXU
NyY4Ie1HvTEUsgr2l/TyqjpYEXGgeo9CbBFuvdvoulzV9t8th4zLcFesXaeN83q2CTqzoLWcKHHZ
bRqFQXutOZ+9uMYmY7zYj4PfXpgN5mgX/7tm4umXaxX65LJCdxnd5ow3ux7PgDA3xpsAiNLm7JmF
Q1AURaTkGVwLIYVh5OQDLG35oNGW9RN1Jar7ZKs+5CxI8S62mXAYQrlb3dnmZyo/JJuCGrgGfYvt
nRuEjE+IgD0dvMHcOgax8CNywobgBpYyTSy/ccng3f1aDOo0qTR9s/sEpwQWmS5qRJQjHXSes6GY
snWhewf0mbJORTjhS+GjLexeBb5PquzMlXsDKM4DWI2iRa3hP8yKSkNw7C20EJfhg4apJs0LHUAv
+IXkmnzRp9DzuRnU1lgJz7RG/aVsANY1X2w7aBR44J7qOFeSWWsaIrNABu5ga9lMe+pnUbnFb+l1
DL6TAWntmkM3sJhuLzS6wQQJNtUHZzJN9YKPNXzp+IFygqy38F911IAK0QP0twvy/FTqy0LKi4sr
Gk2Jt6TKmhAlyYJFzi3icsu2IOQeYrQskLmxlZEZjEYeAlFCB+lNZmbLKQ1E/Tj3UBEfPShT5q9k
P4ckBDP6mF2heUkEt0OZzJe1hMttk462xD3O6gquDK5UQ8p9n82MbswOjfy6ASp/2ynw9CLTVFVJ
GJ4/1csr68FDX3WTVtHqdRTqBkIOtW1+MTZw2TBAz43xUm/nQtnOU73ZXa4TEsXsTvrcoVVhISP1
0xOzT/nGcEv/vuzsKPC+xgXKg4Iy49dPF0B7wtXJor9UQdGY6KtP/syhMJZJYJQhfn5gbocPpAqk
vcnEKhrSBirUUFmiugnDxbfbHaZhy6gj0HzLiNscirp3h9q8lTTmesXoWMy0jtwWN2XB2uqHykbO
za2wgAb8Lf8AqlQNXs8sjcY71MXi9rk6OfnDxoboFyyPqPFdVuzFYKC9l+znZWr09TJ8eML7t9p4
4PxdO8JH7x5GzWV4LrU+HkOLhNcQBTMLN7vQw1gNuQWKI1lBSRdwz2oIRCBdm/QjwfLdLjUCu+yB
vojq85Op5tgjer/NB01KNNCtJgd+zgQlvsDzTyyjLcm35ZXoa5rSbbzq/+ZVAB0E8Yxn6z8MIGUq
62WN1UTewTnp0+n84otJE8tOLXEYtPwyO7bjjUQPFzMGErdZNDc0VcjXSIbSt8CsHTPcDQvbh3pT
v+X1wKCM6XIf8ClZ6Ze6LYfEZuVctgln7KPzScSJW6hBDT6NrGPKunN3c+yMwFZ//QZm1gkZmtdk
KjFEFIekiSeX4mmHWd13ixEukcf8BvrDCIsGbgOVVHj2DjVgkm4moubjx5tPQhbvS//lrfmT2IbI
8joExoWIE2NnWQkBq9y/8Lh9D4uf0TBlu/TdbIxm/kx7WMNPSplxtJKqtk4WGInOQpZUmxffoBtR
SF809RstrAhZB25vtewHPaEjm2xrkkzTNmeVzo9sS35q4aiL3vJZT2tSQUZW27kjpg4MyFdAmjH+
Py9+EWHDe2nsNdmPSl5KLrK6cy+v00SLzdUbgqd0/baFH9ATC/EdLUMYtC7i5jj/fXpSzpsHF72N
L9TnsgmRTXEQ4GJQmncXuOE0jUscFVpL3bbKh8gFOVtpxleVNoTgnicMuTNYgCI9JOxJY2SsVYMJ
VJsYzlhafMGq7PoC+cBmV/Od/9KdBS8UUit6FckxeIL+goODcySArKEPfmn2MFud4uMaQ9vEsyf3
3hZ7OOa97WEWVl+tBxMyOdI7Egm4/oEsyaOLKmqVavSYCBlEl0WIploYdh7cQjwz6+phCmTE6noL
cJ7QvrIqrUyWKP0VmUUVcNge7mUZ7/Z4WCVstSwvPTOQVw3SIvk+gyfbVdFq4HHZW7H6F6rECrxR
lG3Vm4QKmXJMmpHAj+LLmoyvH0Lz4jDZJsb5+omGDAXUbkKlfjeApfVVec64+Kcez8cKwJ2+UJG9
H4FlFsDd1zh31rd+EmG6uqdIZoIB1aOiYsXdF3EKs1ttBUbHNZAvdtdglZd5hd1uuHAqaWCOgMZ3
0VQffIAilwMin/j2sMC9lOpseRqXQWBSRU2czUY11CPcwcUKefJcYZ1tZVRcHeN/CloNzrzxacyy
BeqbeqiV8wBjwqcLmW/Wo/AbpJ523xUp1kIko6mPveIbULEWXyx41/K03WNcmSrflbSjeltV138H
+0G9wpS+iIVdYXSwoxseODtMPauuxUdNVoTwZ2Bdv0rXbYHIPcJZcFPJYMGw0gxSNSZjJ92kpHSR
hNsI3Owu9yzqH34bzgGOInoH1zhtlxdjpuit3CbQ3106r3S091mtCaH+pm0JsGKXN9mekgZPo3Ef
j5HUw2h4pf6kg4bj6ydMbni+lePE7XJhR4wQ2w3pRxjEZmB6Xrvq7IqNNP/mMMTqgPGR/+AC7MW+
cIGS6z46VXVcPh5D8BMMgvDsf6kXLvrkaRDmZE8WHP3DyeHat/0xm6KJeyMhIP+mCy7VT9v5xlFI
76pE7/NTjAxY/GGouiIqKK96vG4Ym7fTIr6jDDvusQ1GzJP7RsbLlyXUAAu1q+pVBO1QRg1JxXAz
nM1jXYTgVf4NR8I5+NCOFNr+k5cc10kNl1PzQlFCdHXy/6ao9jOMjDGAj58bWlSuxWnC1Al40m3V
ErjATW+v8nZ63lrwFvKPmEkP6D3gD6rkIj+f9/jjF4Y8YgjaPfD9AS7uIUvJv7fN1xDT0q2RJag0
Bcwykt6fd+GacbIzn6kkQT/VH9CWdbJ6xuSVzPwuvKbNHZ7Y9xFiNvywg+1MixaXbvgcpxHyQp1q
Xd1Daqw7dy0B7VYL8bKwz1sLhB/A/vSdfIEiFhMv3g0zakkPhc6fbr9oHVeeIXCtJcppUe0U4CS1
4i09VHwVVgA4D1e4PS25oyWjBNASyIZNOqnnKYfgCWWYT+nscITdBGG+Pr9qrjj/ocjC78Ax2E0f
/vC0UU7reyLS8pUc1yhW8anp2STaUzinff04ASrisO5jJgj+/e6AupTCeFInSebQP7Ie5Vtv0UO7
um0TDqoBdfCpjtrBkzPo3RR1/1IXEwJOrxoUyBRuBnOV64+CTYJlG7wdR8o3Ky2IpbtyslCjMgXI
e+f73fE0xAMvYWCXlrWMdIhntMd/tTDqyxsavXlCJuO8Oax5WLsQ8enYHSBYA2lQMSossdVtDKBn
0y7hKiJRgcdCb1nmSrqBbcOPvf6bxz3QYeLZ4sVmQG+KgRXtgp0bNdOIyde1JbHv5fdN5L/W66tu
FbxMlrkNrAtp7huM3durlKctRqfHwzautjiR5/h5H7qdacTHOpRrHuZZETmPMcLTdq7s52xS6ZAP
zgzf8PylrHO/YlrcBOA6Fbf3CSfi3VLeUwoBLO/EJ3yu1J3EYhlkoVHxR4/PDyd259RZHZ++KJPl
F/rDEn+VXifDhf2+3AgBCbMqZ9PgzwpMfyCXgHFFTMMBtUXTwMIpAFtoNoQztJQS7iLDRnX+Ncf6
Hd8e7+lHmMRc6vZy1xDof/RPAM7uLvVXDcmIRX5V8PWJNHMyXFap2rX3kxISqihOp0wmexrYow7S
0C1rzMOKzhvWJ9QzHdofvtN4lvh83F4EPkDiNC1Ru1fPbFd8n7YFPVg1RK4Sk5xXEqYypxKdkP6R
l/zA8zufBY48JTlD3P2ouUw8Sct+kHIdWikECBc0imvM1194gG8QCV4j8XtMBQgKBoowa9rkEgYg
D3nbuSsjVBHRj738vvhjDnxbeo/ZQ/UssgzaF/T7/UhQ92gNet1WoDViyw247QTGYobRfSKuTh36
Fh3F+4N/b6NpC1HMaGf3MRlTpcv61cgUNBsh4KY39eI/u1Iksk8Mz52W1QO3qpYSBphJB33AdXzy
DeuPCDA7kA7H39aezlj07+KrJZaUDyQ2JUkWuvv+BEQfVr3OW9hP9ttY3WLtikB7Brxujs5seEMM
qhC9HljhGc2Tkd3hiI5yle+91VPypXS+IuXxbi4n9BcQaR+L6LKe+2KJFmLIovTlceHiy8g4wl0l
Nc8jlYu6tuXsp9WNXFx9oq1hDerFSzsM+argZ1flWPqNQyjeVheqNXW/3D2ZQw/1OXiGpCyWN+ig
ludFD9t1jyGf4PhynRSUmJQ/6dVODnCv1JPepjFznciG27bCf+1mFi1pnQw3Q0S+nnDYXQyc9dDc
hA75dSQ9eZUQzQ9n+lf5StK8578c4TgICAfigQZHIFQV5/T2GDniFaYR5HmnyQUgv6Dojk5pRo6E
at7hgzH6Mgb0JexXfi/Xnx1rtwKDwrPr8B9Im71CpVrKPaB1rcF7csGoUDjcYJ64sJ+LYTtnJfGO
/KrdkVmOYgsSTAhh4AQOc+mukS4Ct4k+1nRjiAMEz02HDe4Uf1VVYqoMCjgLc757kFwKCrFhL3rW
BKg/w9dqjErctCpiIkmNeFgiNraa4NcXzl0C3OqJTVQ+9Dra5pIwikkW31VNfLQJQ6FgIUdpETmD
YxXZGhKvy49dFlC4JMFHnwO3Pzqd+lkG0PBksXTilIRt1DfaqfYULpBuRrFXD+vG2eCYNCYYGPHl
ziUM9z7ffPWXX/k8IEt252LNEKV1+mpS6vtMixxveJJnFn6fkP84SXwSi1v/1Zc3bz5fWt+NFqhG
5R039fUhsiMMMGGNXyZZwPKI+aUjbLvCNImJEHKenPtLQlV6fO4v2M8iPsGDVCcbhkf9tFQSwqHv
9vGTIA/JUlrdE5ppYrasfEoofhsSxJR3UW7Tjh8jhWpSGDiHZc1uDWmL4y5/bnRY4mlEmPW7VXnp
WL6o6aGgwtRyJJhbXDPTHIp4Bd7HOAzTpoaNC6YcroLLF+c/6p0ZWiNSy5I58G9HcZTmBwbOwEFB
YDQ6QcMpH3NYJQBdvIso2veDVXFtgeWpBsXZ92DdL6YMckHA5i1g5Sf8u06B68dulbzyZewHW7cN
Khp2pedQU6WitZmLx3iduaYrL50HwgP64j6nabEQN7aMXwHI/s3F/4aGF7UrsNxsr7h3GdWmD2Q6
AQkfLpLb8M+xglBbGEupK0kocuOWoF7ksMkuU11Rnfm5eVUDxra4ZxLFKTsoXw6Bxkia/imqVb6l
6G0ILmj5R0MuXapvWY7u71QvLhchaPsxncWbRfrIWPmwfeGODm70uevAwQJpf4cWaFUJeDRDDiVc
BGGwNrV8Zm0BdtZNoKmiJiuveqWmKxxFRVWrDut9v4PAiBeHNKtSYH/2d3dFLVUqQfF+3JKWsC2a
mDsDIK14k9hdn7L6iyI5Nwvmfzi1XEcTpnSYc1tqlm0tVH8xE9vZxMCJkyMGX6i6RsWnJmGm9RuM
MYA+LWsejTSOazzZ+ZMb4Awn55eYZdYN0ATvX/pi9KtqmTvkzkV7rOvipxbvgUCufguGG8b38LUf
sBCqMUjmlXzW8I7LYOm63zdaaxG/WnRTnY6j3ch7O7c1eHixo5FXxMa4pdtpkpIK6JKUIUPum/kd
8vyltckZSu3M7ujSinwOzCZFlma2RKB7WukfE5UBAeT5nxiz0HjVXJHFDmhu25d0wVcwWArUXCqg
q7oKKqiPPR19BKYBxIwiUmHT7QM1kYDV+cUA00R8c2dQ6xWdUlQoJDMPPQrf2wIpoIhjxsMJOXg4
yhPb8DC9jbsNiwSQihT50K/x5rmrJgorih44rGi3eLiY6P6ZLWX6OCXCATwsmKfnWtoZJTKTQ8hn
PqNz7tLY6TcDjrczcIoNlv8BsocUs3YIRkeOAsdVGyxIOIodZLtsXfb+MW6IWC98DaJRlU/9I31x
cOu+D+iqpUaondOOvO2gfX2bflGqiJE25/8CtHTB+LSzOFshesNjGWuDNcBbepvhbqyqkaTdSmCX
0dAvQ7K5pt70zthWwA23IyWVm6nMCq9FsHOu0WVJJiAXwUtmEY1XkxQ/3Y97H7B5kxAtuCum8xL+
wfyxRQxfZgj4OYtw9+zokdYj3um6IHjoMv4doXEvhcQG8ATxXjVVYtjHyTN5HNmA2wrHIa95++1H
r4nj9nyRe+jqau8nozedvj/031BXrc5+SF+C1+usZHfj3uCFC5/D6GbzJ8WaGP8kqTS4c9/w0OfQ
7xKCfh9rlwDeoTa7QkHH1bFwM5aIrCRNEcVdsxQFd5OeF5QOOSwQ12MCOGLTLeSUyzzTfELqu/lb
kbyxmrSi2BpX64I/nnDnLPp9dCeiCB5Hs16CrOjeetWamWgmfUTdJ724loUpykRuTgqUoCnoGIsm
rphBE/drkaWWzTn0AwLtg3WCQ0OGwMxlvMehdQNgvsxQ+tHR6BOiwxgbVIYo4UJ+ti5GMpZIpXUE
G1jfwdYd8ofto/rU4Ao2o/GWPPI+r/XJcWT8XvzIblyxU22goiCG7ughEOJG7zoGL+/Onli/oY6n
BQnMLvXG2vCYe9ZZ3B/nDdEw2zlfZ/dWRM247SLf/c/MKhs3I3K6I3Ga6KvOgp5AEla6rkaVHdkJ
MdW4+uOpqg356MWZ8nrgY0dFZscxiHm8kfYpIzHvpvgT9mYby9Uy2KkeGQK27jG15LEh4jc/tXMl
+/h+EyLEO2QH6EW8KGX9LPwNfta7rzD2MW4an6HxXFqzjIL/q3eip9yozWXif3AoZNKTtkvnAYTj
kP2UFslzn2oa4hwlEjEAdD0g/YfQYt9e+JkZZJOMh1RENU2YTwcMManUWEIOHUCzqQaUPxVtiSVZ
ZlyBJX1V5n9qowFKd35clLqle2Z0I4NJ6s4j8WhcBeaFFGpQDOdGSFJtxp2uoX5txwO2qeQVygYy
G+typIBz0PLfMYrMvzCg68AmP35G9S2TQdWNOJ/PqhR4nPOZVm15V3CfxykhEpDiNxATRXFqQH3r
kvG7xMWjdhA1YnZ95REhZbWicalVK6siu+DDzngjJ4KRdp3G9fnIVJiFhczHeP6xhFrniIzlgKPu
CwRKDVM9BGMegQDhqwMZWMyYGQK4p+Ed0BkNBnSX7LVoBD/9WWnI8uh1Cib/RnYP7QAsvc/KO10i
g0fjpvPK0vBdtZywcrB99Clc9NQSgKxbRSdDqCPxNEtCw7kF7b47K4uCoDUw9U/lYAb3TwspUTvE
PH2VaWI/nEDE5G9aftJWLf/zPINx32AVA5mu+OOwmEh5LJuvW4jtT3Mwt/t291N2vdV6scjfqdZz
cAEMMgzMaNAWtdv56ckX/zIRZA3Z0A5EKYFpsWFh/db8xXFGwPTEldyvl2jro/jSU4xKUoTLFoOT
Y4wVx+YSMfqpgJQQBOoLGJazfU9QwAspAd7KRzMqBA3dAK1qMiq/RbyWWfjSeMQjk9QY9a8AyeFE
rZ8sfcWcn47FadWlURFsk0259c8g1KLFWx6GUAvJVsxWIpFnGgosxwbHOj8T/ZA23BW4MJ6ubcFD
qX79Ibtkzsa7v7MQoy/zL2DI+BPIahzjAYxewBZf62bFs+uEaMALTE3RwJy9CsLDFSC19bGOZhxA
4OM/sT17k+BNvzpvp2zpNyPUTWYmjKw6X/kkjYYT5qJL5CcLiyMECrYmvXGJojOaqO5Wtvy/kNpR
zt2/w0EcGqmjGEb25lSHeCnRRI+DB5rDiiX2lwMYKkvQyTbinp/tEzPW0H4zN7sOMZxAV+gbuHWL
bLjBKbHAByMJSkppciUp55WREH4vFT10D7MwdWzFexWx1dX47cIChjnxqO9WL/0QGdl+b7E4/PDc
Ly2YZrB08VgWf44lgN4IeKG3MP1l9M6QLBcAqfY749wnoNpZzkM8E9YQFvKvZK8wb46WTQHRmMLs
qd8k2owcD9HzSxpJjS4pj+4wjYCheZPIwCdKzUnnuZUWoQrVqRasRZmbS113MK3lqi8iQzpAs2LW
2+inzi86jmlHpeROMxT6vkh1vJ7zScByXG0VX5X/KZz3eIBvLpwFtDdo/jd9sMJNuiGg/oP8H++t
YKq8ZWHfPYxuy9nAFhU6yzDsEKLyl7csxbwv2Atpy20tvYZWeTwBajXEzpCDCo7ZwnwpR8l84P1S
/x0EzOS6we1KSC4FfdIp/Q8Z52mg1bEJNeDaMhGjlXTYJAEmSqmARpuKRJXiKuxBDa4be+HhbtUs
PRODdG3rr5nfNeEA3veeOIKB0L+sGPJ1Qx3fQkpDkNFIZmtlAmpwKoa7n58jI/q69Ig6bdxAjqYp
Mn0TUPXA7iRgf1bTiZIXqKog/1vYYPFVzxpuhURkcOzNMxaGuvxCHvaWDwI6PSOiElQXivpZQGh2
nqsmnLZqlw+vKsT6G21m8tyXH6kUm2SYJgZlvtxGqs7BKueWksaW8yf/z2ORiZN+eGn8cvtb3RYe
t7Vl6KehyT5Twwq5WW15ZW2gCzXHv/nCOIFMkP+8N4XSpA7sQ5e4uQCAk69ni8gFMCQXUofbzn2u
j84q4nE8caH2XB2nFg2pW7znx5nkobN6mkaJrv9fsTVsG4UTtvMo88J1g17FMFSmBZpY6bhv+dbC
rhjGETDvotZObTGuePvB/nYC9bs0n4dSVTZlgaqnPGhM4mOeHE+jBqlWAYTDsFMiOwQ1hLM/XrY2
p9gGrVyENarjGoILGI1S8vN7fS6kBwUinYv1oaaO3o7C3qVo8lRNeGQXB1WyqhBnJY8KJwWn/0/H
4Kh/ZnnfCx1ijjKcu/coF0YtzuTJN1qkMGjN9VNDYSm+GlwbOcc4FFP8W6EZ3sqkSw4FmPKRSsUy
QqPXrMsZ2esvDIUKEw1Qp9W0JG7M6pvinKedMJ+uFFJZBa/OiufYLQKXeDqCwgUQl3eVwOxq7g6R
0sGAL+mM4WX50yztL0L6NUMuPIXGoQaiWSqGUg3ivcQ3jVkHibZib+sps0+uoIV+DN/94VU9q4Bl
M0NojQkdiNeIH6F+RgM31agKJMIM3ZpWo6/tgwDWslRXt+ebUTEBxnV16tQIHFzuV9R60D92LMXg
GFxnGQJ+HrTeoisUFwOIdkfw6yBgeTtyChDEXEFm/timb47fihMNVHXT0VmXo0MsOSnTuHdh5QIX
fIopiKCIo5A+PoFHaYEPiZswyCJMh3+aTO8FyohSAZ4SGPvnmQE7MFM4YpCrO3EHTFn8NCCLk46Y
FFYzKYc43ZAnRVe+jzjwjvNgWoSfB1KdNO2h54cpl8wuBkuvNZEKqeB5AzmJ9biz6JvSnxfQJc7f
ZVsX84s8imnJVm6s61YryXKemzkw6jgbP4QY4IqO/JDWOthRhO2nHBt17MkFwUupmNqDGZPOVd2D
KRSZTN7Znp+YT/yws8gJkkQl52lXOr9ET58wBQxfr03n+GvB8LEinPW5gv7TfbyyEb6Fh2ZsQmxh
TJGwk7UCFvVTkr7lr4vX4fUtURERHEWUK0+jKMiWXRROEtJZXNJ3OlaLAZYFS/t+KKRs7NQkJlcE
hhP79A61mVOmfpr15pklSz+oU6u2XmjnFYxPXzTtHJ6qSihlgdUo5JsngTpvNpor9/5vqppJk25I
/AtATByo+atkKdexJY3mx6BfJSYZwBjJCTujd18RMAreOhNgSvKun109gkHoyI6gNEnympEFuuAa
v13GsPzG3hWozf9SToDOEEWX1/z7CtLxdmFWufM+E6QCN6W0to7rTGCk/p4zm6fnXAO0yMtKpY0y
sj3A7I5uSNDqr7TxorET1Og9po8ItmV9z8zo7aEkJg1wYlJptf9tP5lGAHv8MPsU8BPo5L60ypdL
6CfZrdzb+AvAXipsjBG9HOGa/OgeOx/HRh9IB9NSmB4IHwvPTuBT5ZhDPF6C81ElQY7R86ehiANm
YIklBuXNuQ2cYdpXoIomxGJIYoRr5BbRUIeINJ2L2ywWP4cLypYsTa/Abkz3bvVAJ8dGC//2axk4
BZBlfRn7Z05vagfHaxs7IlBhYubIAhvqOVvoMd+Q0NrU7fSD1gCd2Ms34eGQRyACc+rDk5vGeiGQ
kssBkQkzT+yy7VlPu3AZT4P8VSKYrtLcfDC8Jfo1V4aSlt1jOQwVIsGRxVLLnDvqeXBINkdo5ZDX
+l2lK3L5qZyRkmXyFRUPHvTO9yBVJ65LqS0deaL28RdO8Jf7BGbDPP7OVSSlaNWeykCYB68z4hpq
rUFbcWPcaVaA9EEPuE/EKm4jHDBNbbFhlZRVhbPa0kQ971gDAPM4uTClOLmb/e+9z75zLoL2zSNm
dlAa2uYgizDDP2z66ENfBT8C/i4yDIk75FxiUJGeeVXXKcoNs1xbKhhVrk2NkOSSe5JSRWmbqYDd
lTo0ZrONubFd3d1HtQbrq/Y7UQMVolJxhhcp/trmDMkXiDxEmf8eLmmtvAXF9N3BmsGuEg3tKimx
LBZrmr+GmI356CtQt+nKL1tMeZpNeEiPBNMUDe0PeOWHm8qaX1Ir50uujwqsz3S0IyJ4mVJEU32G
R6TpDV1z013/p43lhak0KzZzdcn9yuTZDgz9Ka/jUwPNxFST2BxnH+FuMG9vNf3Ay9khlzuUIDH2
ybOuLiSK0Wc2I9tRsljM5CVluRIkSyFdb02bq1OhsNGVile5zBrRTxKjwPzzCTmenqhUoO9cyOpZ
2YqXuwi8VraKI+SFfovFchS/f6tiC2D2qmnrFoJ/BmeJ/Nj5ReH6/2pJyQxY4N7hre8dmcC2zHZc
iWfB9zekAvXQPBltFSVPoaLKb0FJVcNxv2EIi4bHh/+N4Hv83CzxzA3ZbH0bhJJpUxxO9kZzCTF1
b9V20CVOyA6APYVByEUjwvWH/lb4Gj4rDWU4KKTPn++eOhpYTRUdyXpk2W0Cw1F95bxb+dx3A41f
oGZpqRBQkHVk9i3vXvSNIg6nbvYeikOjgq1fiINglajf/Usjm5LRYAMBzQ1p6w36Mln0Qh+eGemD
77iaa5hqns9UXnZDFhANWpL7G4eCz5fYGOITBa+p5BIrCPgtVOkzTM7l5cjwDDsw6r10YPJS/Ice
yDZoqYzPKNBLK8EPlXTtqgCHpbJSfZew9UyPrwTjf8u1kFunsYjUgg9Eq5BiGMmNHkLuRL5BFSq4
1MjDWM4C7zSE2vI4cKdhRCYiSubkrBOA0VJhG7IIiRUg8J5FPl6aIX204/kRu1ZU+ctR7Axn4ObJ
n4fC+ClmdSFuk5PKwxt1JvnusiL4eHIeYbMGhh5aeu2HwfxZ81/QnPMyMa851U8E3wAg3PdPAFzo
IFWSFp+q2GDZ2M4ki81uLz1Rw+MyBc7NlpjngT0Hiu09docl/ous6Kpb5hrJk+bTIT6rvPjj/zy6
+5nvlGaSXzkj9wU/ptT83KLfLgKXBllSrdLu/dj/vctIZkcjrNZOvMRhyhzKbDoS/0a88fzRLOcE
YN1+tPcRshzkNL4lhU7omEYdyAEpLaaYwAxN06vLqHJ0rTCY/MEgR6Js2RuLmZtU2UJsb+GDPj/K
LuaMLghVMxZfP2efvTNZkSbb/VXOox5WKxg0L5wRv8IUzw5I/7RNbE2fBCt4yxGBqePGoxxrufLz
AeIv1H/Z3v3Tlr27cpMy4X5JQ8GObEym+Kt/YkKyEQifojn8I6SuJPi8Nnyu9Cs8UBT2iYtbi8Z/
/VqIzxbWzhyLRUSnch+T0qntc8c41ToGCYDHCBbd7WTEyP7Pb0G5EJrTqgOHphvGetIrNRHN1ioh
sRugSJYKtPmTdNo2ZSoGjVIskKkz7gnE+T23uFJjle3y/WUyvYTGrXGtBKOOyJ19NbSvRIsABpXs
hwK9+9h352wYsPOmh6EvMpq+3AZf92QDXZywN86NHmOnzhQadsD3tvGcefmEnNVYUGs07RJW/Esb
bAJkYaiIGDlFCld4/ig515ZrUy4/jtIRX1zwZSBm50c/2HxwV0fYlyXVBz5W2z98fz17rLgLm94p
VVPGh8gpUhaJw32q8xMeKEM77oe55kEra4sAFCeua3IYiaH6CwjDZLCwcLI5OoER1UXR0fJb89Bm
OrK1cBOAu59V9gO5oMnl9T1ZlNzWuwz0dhhDz6KCJ21JW5NpcXGlibZeY0/33f/sAuOjig0gB1EE
3Dvwb4qqi2QZuBXpDd6nh06sy2vQD07p5X/21In/dGcsVJGfsvBqkNhTK/XCEtRBHVqWA47DCsvP
gCmh+5CbGVXHnpV9cHgQA4M/tapXy8JKMoLZ8Ou2AYQIhXFPwbqstVsAqFt4Ok8cEeLe3E04idzz
DORk2QK2DYUscI6IIkUAPnD/FVvTnsBDVW0+f/HMepEP0MUiNklmIKYRuS/EpAhl6xPWPHxGqIh6
Eo0SuxffA3zl4HeckxgclrbcLuRAlJphYbrOYk6EBre1Vkm6h2YQv7rDrUTaciHWJYgw6toHIFC8
PCQpDMFCpftvZ5bnhPJ349GQ2P04jy9d77Nq7/5iSqLelWw9Awx6YBHLNxdfmR1oMIfEHRHQQkeD
Kc9qbZKt5IovBDJOEhVuFxEf3qrppIbqFeQPV2gBQFNFb67pAHGpPb5Yd7JPe0dURTRsxxVPR6bd
Ktu1ZMNF3wGPck4vptzi9hL3UDnRunDhrykyM+EQwA8RTSn6MmWdEU/teke6NPKhkz7anaSphI4y
DSPTzqU2fboULnhiwPhYsDRpY4aHIqK+lJMaOxzIyMNs/gYPPMTjULpiQW/ZGo/3W8hAT7ArSvXw
CtaMNpiNl0tuLlnLYX5ocOSN7U6/4cu9oIqADEK2J0qyYp9JWwCuj3DMXRwBMWLyeuD1SK0qKiDL
c4XXPPMMIshXru8D4bUOZbujgj8CspGiD4lyBkmpVtOYdV73sUYLgZVpXJ/iVC6LKk4jQHNMhUl6
3Tbh8cO0apOEd592nVFxk8fzVEsvql4JbtnYYSeHmRNuKsyQQgH/Df5FGGIiaTukswmfEXoOD+3w
5+stNRFj5iMg2VKSnkGjMLHsJYG43aw6o+eJNr92AQGU0twc0yW2WzPp/pSyV7G8XKUs4TwnagMC
ZFh8GULjPEADokbFIQpRK1GusVwYwrV9657rM4gqrFvDFn8gEiTsmeQbrkNLXuLBSAolVfHAbSX+
ZXA+prO1KnCA4Evq5tgk1S4weyiieIs4LNdHRsc1RTWQaMByb6W/PdyUnbwgZnuplij8RJw9lzUT
yTz7G3BZPoikL8/fvNz9uc1pNyDhfMDufWcA/jBfqC0d8rtVSvI84qcEe2NEMUgUQmR+fS28Di9u
brd0qPvTCEs4VXmmVwu/MksVOb6H6SXH37lQExfm0/MoC1p7YvwrIrvOVb6RIBb2M0lF4y+HXnWI
6Q9Xlj3M/Z0mm5pOEnKje82SZQVDNHU1ULaXachElIpRmF0mD6Vh0fqSgBsr4IMERwBdQ7DXLzKW
mIx8UDqzkzVT4Ll8CVCeZ+xfGHcnAt+z6HnlhuRVXRSDUKdmbG50jhSsnEI7EL4j3/6NqPalR32G
V8vwVU8N7Q2FjLMVhrsmAxJCgrgXtVXHsr1lVnNadNSnE6/ky6cy7iW5NPowRTPi84oGOyJnyR5R
mp0zEmWigbzI1NQHEq/s7dHMDnSNjTS0zF/H2e54yYy5//cL4qExzLHt4WZ71vW52LLvjY4h1b7a
tbVmbGEdEF4iqsUtR9wwYqDteTZVUH9knBP65VcD98UvyfDgBvriXLybYlAeYc6Rr2/u+E5rfDUm
j9YYKG/95XuHE8UEaV2QKlixMNFAfrSYfoMH482yJVTgKOBsvJ4vCCz6qu4uE3iWa122c8E/1Dho
973Inde7u3H9kmUnxcokuXZuSdZJlF/7e8WBiWRgqxs1fSB36P3umPoWPIpUkleOpR5fy1wbmAMD
af+hIPkPHJmhVTddg0BysCa8Qurfv2NU4Cxgs/E0INLiAZ4Fv95EAA0dMPr1WW6QH9+9ukS0uk7C
6SXUhZzpo91erMIz/J314Y5L6UdGKM4vOd6A44yUij+xwP8Jqmx7DdODb9kfteMX7J8FgJfmhAcE
hJAs1USRK2LxPTtOF3VNLMvYEHo/8YyAetqOQXckyZ3xcLD8MQTT165pYMNYkv54B5NCkI6blGaw
qcqE99WrUAvoxgXE3M3B8+FGNWgnq7m0YZ01VCq5DzjDVMXJ9IKe6e3T6eQfRISlay2W0tu+n0Np
Q/DyWCIWNBvv6t3GC00f7a4CV9qgAp4qfH3P2iU3U3Oi+oNM/mRday/T10X6pWhpodX7UizKSSNm
1is4Bh+zNvSMQi1q/aRU7phUXVWSBXOoVAdpUB2R7J6REH2r0S6y3zKhIIkCsEDj/AkwCDNqEcPR
Oa3nl03XernFR0g4klOn10Nd62PSlJaGItVB4UdJ1KiOu19eI03b6M9/8cg5sQRjkaiKk8UdrI2Q
IwLC1jBbtkN2g7O30ITuKDCHVLpBwfiTG6do0r3QdHe19GxIIMNRf2tGoKkUtqx9oZFR+esi9cKZ
BJCDv2drikX+u+t1f1pr80Un9uVNQfT9qvnbBFa/pKAcknzNdId74arHp1S+HhUlBpNUk5rHEpcd
J2Z1dtbv7VDwafSWP0pg6D6OmjWfx9A3yjdIu19tZYMWwYeL9f+nLOtW2HLS1aFTnzOa+OQm6J7C
zmgwwAAP+Io/zw6sJ5mMucvDuCggEFaDP8QWfWHuewV8ntjqp2Aj60Ou9HX4nMeAkI8Qh8Cnvzhx
fzS5ccHxk5ozZkUubSZ9N+J5cU/UJRc/MTpFPv7GKZSDg2KNsNFqqCZz0gKtvw5J2LQ39Q76dFyM
mWwiBEIABxvakyTiOWXEVNMIPzQTMjBVTolNC8R4O1X0VKzhR7L2DxZ+kTfIHlL4rXQ2EMmctdGP
9yiWOP86H7LUEbCNCf4xSf/qQFJKO3rmHddYTvlHMBeWTpMpgFazcROruvznKZQTqNjOTQfREw06
0Z9BgYWPRmc+8Ti2E3Tqk9WZmBke2qVSo32pK0daaJQFT5H1uoy2nTvnl9wvgq4LrhWsC4HD9TFu
YxxacEIa5Xk/ryqadHjjYHV89PZvHFgEkxURvhJEVbliGbgUKCKAWy26Fz5B5UJKJp7E476KgzZJ
bF8332xuMRACOhg8qO9rhA0zNSkMhHIF+DAd43ezexabOQCjFGCLJaoBz7MQA3iFfmkVLtz9APNk
Y5sci5YWFPV3fIMVytlPFurjoSfL5F8pRzE/1y+mRB+2ha4REkvqRcoqISKs3SGyZyY65lb+hLOl
8rlX/VBHf4BE9eFjuiMsFo9SdUj/i8CZx2qBYdhpcsyETZQJyBfgJb7QjGQHxV2tp2tHj11hfyzn
mBdwkqhICaHp57M5nTazqkkDpvdGzIjteQfrk45+OE3mrEb0PtB1S7xRicAke9MHGl/bDytelFiK
j8DCG5I98idpKAZoX3PMnAeZEOIWikSnTrXnPbP0OUiLabnsjrxOJ5bi3u2X7L2L5gJmyEmRDVvw
JG7w7MnAe4Tg/116D/+TvNCJBToKdWhRfbg33osy6NvChyIS373CEga1LaOAF8Yl4XvA4vQUNJsY
2AiSt1+yV6cgpiRJz3VSHiJx884V/MaetgO6mhqbo7XJrGEKPgzluNOD/HzMHWukvDv0wD2WHRn1
LLuTxgAwVFkobUS/OE/1idSL6cRkyYoiDXRs0KEM3pjUTsgHZDTyT1RT2760ASQdWfpYyw89UxMB
fgcVNYzkfvyH42BlZaZNlkaI1KZdsJs5hI9KkXyISQfBcZNezdqj4w+hqxg9iLtTWz9ACWgNyEAm
IL3Ddo6Ou/3Z4RcVPsrKB2oquMD+zL/fvkdrPjr40cOKKQQHU6lJVHAV3bAwlnSP0KvraPY+7x7p
C777u8bLlywCl7p2ExFP+NRl+7hMPK1ORhw//u2hoCyqDE/LwY2llSC8bBMntQ+sHLA/unUcRAW3
tS7Lf61CdGGN43dRA8RbwMIRPdJNRpmvzIa2CtD9ssVDdjBvumvKKiT/MQBc7TmHf7XpbtMUJwtd
7bCGkPq6FJ/s1tp2rIn1fb5TjE6UMZE32EkdDsNTwvKMbirBp7iHT8Itxc4ZO/4LHyFoJ+QjE56h
MG6744uQdrG96vzYBxETuOrZlN695imXc9py7cvruENetYXKk9zM4eI3sgB/5LZSaBTJW5lQCrop
tHVrS04FIp/U7lhf3J79lDKROO2hzUY6GDx+rDHJscQcHqDlng5Yfy3pmXib3M1K3ptoZmjfmMvJ
JSLyJdylsvi66Xb9lFTbmJH7myrvqPATYu8kCCy7KyL7jVtEZiSSDv4fe8wKENAujP8bkd4bYpSi
vrpuCkgNNbZbH92wsBIg2mlZd0FWN6G/BgsVIMk5IB6ExUY5LD6ill4h9Zj+r5TGD1yfGcujQ68i
62ibC/KKt+qC5shk/83wZ2t5j+PihuT0dqFExfhYHjRDAUDX6X4ZLlqyVGagW8E2y74Fo8bMJmXJ
M7orClGxjXWTZ8hxNAJp2ZA2X/btNRjYs9CH+vFrZkLnUsBjqJcH0IMVLDf3EQGcVChu4PJLTmy9
DJF1AMMpSQ73K8T13iNlXecmm+v78MMYkXpKYDG9kQgdu1A8NkQjbtHpeS92RcuyWUujk1iNpvkg
2a0qZq2b8rSWt+TRTTDJmReqcBMowkX6JJNlumGNncEHr1i9WK7YQtoHFJpMjP/Wpfjt+qc8HYbC
YQKvfdrb/yCpQUbTNXwjz8DAlQFSgBFyuEGvZQisuMqr/TYafD7bmafzapEyKlzoHVU5HE9zDPxx
2PTVwac2rjmqk06lHhShXAgqpUztcLk0yQ7NahJ8/2/B1BmFfVjYYF+13IamUas9S7g1feIr+TKg
ZlORgxMi+mCmqM2l6MtjVNw1tcvZlw07p8hpTmZBsAUEUPiumIFyFyNZMRM3o+8UZvkylbac5GNp
f+FqkXdq2ukEfZUYZYbRhp264Tp14D5room/l7tZcpcvjAxySKGaZTr/rlT6YKISIUQLWpdDsxnA
OLWZtx5VjoG73zW9Qthq+su5K/pjyAgjvkvM+lAf/O7qBkJ0VWJECwY48yWYUSfv/9U2EtBgxf1v
+y8x+i6vWfUNsj7d0QwdV+lswMTHFfBnNZC4mmz8LE8LPhHnNUlVJDO+2ICN1OBZoBy1HBf/vV1+
Ru+OBF84bdsXdrYlhxsUzpHNgyEZhP4co7ho7dXZH+LYU8D3rExiLttdNfJGYOB7P79mWnE4Fgc8
n8iR7fMOwCwtcC5SPNjnlG2LETaAMUKMvZfrhq5i591OcSHegaB9ae3SQjVdDTcCfVZiwmacDNvJ
kQtYkTFwHEJGDPKfmBoWnsqfFXodbEPvUume0vyBmMnzujKmTnnYD+JFi5LVPYmcUcGniqQO4zoH
UxQFyWhuAdP4v1fns63tSrz6ufBQtcgydId4bLhIsuXtRY56is4Y/r4HZdkOtkF9HMOb3zD2bf2n
FtdKQpN2Je+BA6YNDiTb9C4TevXWpFVELfqk7Bkjh+mi8MPJCINz1jk6mBFPsOFpxWvByzmS7vq/
kKU5Dl9MXo5bknQIAh5vZXG5yKF4GhEJxFkDvTfL9ZwjxTKiq5MzDZL4a8Vb6ab5zUwofw4CxbDa
/MlreaITX9coamm68I5VQsFfeBfQgxKT237WpG4pvSpvpARDp5ni83cff2uXQ1eTe83MlX4atLwp
/Tp/pn7tHgmztxnCz8jumLmJ50Gj0sQ//snCrriMGaeJ7jvPbri7yezET0jBvWu8R1no/3kZ1ekX
ti1WscBgx4+x+wJFeQsHUhbEbHIJvyROVW2uYIY/9gbqS9esCtfumeC5PyvBhf1yKDtwY9md/zKl
bWVrUFiouRgzJAzOzvqRQ+AiVNyiS43JPa5OFpet0Y2qEd5YoZ5vrDne3o7XtxbyYkgmtZF/w4i7
anEFCEIi4d+rEApSF/yR23petIrO0n/jHL8ZBJT5FbKFh4cppNG8SBOYVuvf1jrUC21hPeJVjvXq
lLcBXtF17Sfo7wGv8tFmOyWUb3Kbt4FKTo2K1OHMQCxwzIHohECaXF59kFvrbrYfGRpkoYsQSaam
weRunEtHBNChrlwFwMORAEl4yVqsdvX9DlaYCHnl4tZ2+XPDEPZRuC3eWoBqG3VGpNiH424qO0cG
Z/oaiycFSZwgBDB5oUtWB1C70NhgyIyAwChDw8GAkxqK/yhHarOYP3PoJ3tz8GIHN3+EmB7fzFw9
788ecrZ0vKmJntEA1fOezzrYx+xm82TDvF1lGdqyWirSdQkxtQFaVWNKV8NVkQNynlP3eLEJa58J
RQe+CQQvvN8e5UuDR7ob7mcDyXmK86feertnnX/NrO7NUGNW9DKWCNAcg8O+NgCzaJThwxyT0Jp4
K/28PnNCTt40I1kLAM5bjKy0rqLB8UdbqcwaTlcOuGfJrUxM/aWC397Zsq3newBs9h2BvrjWkKKY
/PvQqrE1ZH0pLErIWp6Mua3/Fuo52UkLRfpUoqF9winC+ceiP4jbvIIhPkKnXQLs1W6pMpHkiBvH
BXCSXxwuV3tzuGUjJI2mJgEL77FiDepNYpQIwdoAGSFa2eSjg85Ay1JDV9WKs0rEjf9T5cqRnGXU
Fgc0c7GH8gUqpka5xrXuDP7mH/EijdSJnTf8X6OHHt1kQJcizeIrN8JqoleWwlYGBzR1MwBq31Br
KgrBUN5rHaE5KQnPbznknxfoPHrMrdHRVd5bt1fnWyKs5lON86dBG0+4p2Vcizm8F1zRgPIUMs28
EDhJHe9lZB2uuwBfNLA+2ErVVQgltjoLdbhN4/yUrsgr/On4ndoxi7bdophcvSWX30phI3XubreN
66hxHWU3NYwrkCFXkFAnC4jBp2+Nhi15cT2y0niFnMADXU7cawi88gQNV4AjV/eIs6uTTqTYu7FY
UCcgnioDFHuMjzAcYtCGcrFv+G6SQyXaxkcB7q7owxSgUIDSwGG5WhLX9L70DXCzXIN6mA4GBPm5
f6Km81sLRLH/HKzRzuvlb3NjS9/uhdgeKpe/5pXRFH93AIDJuT00GAzhale/a+ZccEzP9skP6cLy
zReXJI2iBJOLAuUa8TD1vhC5jK9lyva2P4DnbjF1j5NjMqa5VGXCT/oBRFauZOhkiBQzXhb/5Wrn
oYrjFKUaBUHoNjVpjzX3RvWJ1gfftI2dDLZe2PRf4fQ38UrzrAU8BU7yzhZ5/yoWYmyPQeuPdRva
ZTBj1aBi/0OS4f0pGeFmEnD1J6TMFOfTNs8pK2Sa6oFOyRYt4cYtEUXQ5g/PK2Qp7bBf+YrqmxrE
AyrISBC6+Ya5kFW2uCY7W5YDdn0arwCPuAJdi/O2l41gs6EdD1oVFIkkrwx+bPk3sIWdOuiJg79e
4NifPWQmpoT94IqwQ+Uh0SGE4Ap/+G7KXJQllwfsSuX0gXPYOvM2j7Q7GWnBe10A2VHVqgBPsyTC
68/dpL/EK03DYoAbMv8qunxsd2VNiEGq9/T7Hsdq8bqtdXXiR33lj44B3zJNk1DEKoTEMLiDY4EA
gzOw+3mzR9wm5cbm35WgWA/R/YOipPLtAQHu7IebCgtL9o/pxwWRxSE/GNiGWXlmLqfrpqgi/0O2
VaPy5jODb6UpZ6cKr60Sj7BzM5HaS6JdhwTWc2Jm4p+Xn+mzM6OgXDfzIu5BIs9qG/ZptnjMATSG
/qoLj0BJul6fYLrU5QhQk+fFRNhprw4WWm8KRbNSTFpI9UnBmj2ixx3UCLs0C5kYuiybhoWhQl2i
na2KkwHGVIDeo/6hmRjxXFwqmIIlGe1CVx9ggdOizfimQmtP5CH8/cXOsxTDeWTRWbS600gWWj5b
M53i1cliw64kS/qwY1VABgUqC+ymQXVtULxGMKP8gXdFKmb/UQ36IZmjIPm1djbuba3pGnyuVRvr
kYQ20OOO8SJzkybMBoMp5FkC2LSVgHWYTI4plyE8Pj0WgFA69TW3Myq6R11rv0ZoGa/AmKQ3o06Z
yRZpYkSLpvBElTCHybttFvC5g1IezxqPxtC4637M4LjpAiTHOHweqPH3Is9I55J56kDr2FfE4grM
crOaEsFokX2qJAm/iY78mpoAP5TTfH5ZgJChvhH1zHV9+RO9BmTgdnSKz3Aei9CIrVvTjfUUfVhX
HI0VcJTfFgbEf7A1MOqgfceTakyc7SqYv+Y+qoQATjPheCO7MhnaF6uBy4Of+pEGdP6cTtXlNNeD
WefJ2Mv9sXICNDnepEfDocxzL8tSvG3ZyXEFv2ViAsq5o33NHH5h+dfCZyBdy2MUoMhhWzZ99H8k
xizsToijQMqg0yOEP6sN67/wtdzy3ZFDzjNiudIeNv8OOzcARrMmSpc9yZ3BLMK19I1a6654V732
n9P7uvYJ7D2VIRP/uFGXTL28C8lTY6F5TELaYB+ToYftxrGWYAaWORhR1QjYUloXsiaguLgdD6XY
/j/Slb866BTdWbezv4IUl+f4br5gSwZ02HFHdPeVs8SwTQtb/yHfu34SYYKmTn/63PWhfpjBJyax
UlUAkpqjWk5V+4xgdEK4tLNBxB9J5QEN5TQNTx/yAy5sNGFr5DSnofc8MdawNma51CzpjgRnxFYs
3b+XzEpDZjMBsL37qoxO47WXsCnhLxpVaYI03ptUnY5F0REKBXgvkHUntJXySKP27a0TyiKgTMcQ
avBZN/N6/ukuAWVu20iAs8RBM31N07ni7KV8nBq6EBxpAqoCfV52umW0byHa+UvVqTobIQdIO7go
vQHB5EWAjziyRD7tcBugc5jDTxyOZKvMzGF3Y/IfAI40+nE2n1RWrtWMc3tK96c4Nt3lmcX3XYP2
PVm0jeKbQws6V6+FSqvc0d5a8PGMih0xd4t+jYJ+6CcQ8kSaWBJOmW355xLfhGmysAehNjILaC7F
SDGKqY9Q6YtPmCZ9AdX8Zt6uDX6jqRnv+E+MTldCXdj7K8HDwj6Cn3Twquosnq/6vzJfCSSbhTjY
OQ9GhB4aaMCDY9iJxD1Q8ZML3+MI/wuzwmHjTMGP3Cz/7g/py0NmIvnvVbptiIORcm89YyBx8cVf
ljljb4xqHqVxcvPjfj5L9mvn692hzAilqukzqdAP1QBheNXnTQvFc0q76xKSAOcCKskWpGdJDE55
7t4g2pbjS317ZOnz0edHCX/n1UT9Bkom3OMXHXqVqDsxZthpOtYuIZtrhMqELeawipx+TwgTWsIu
wnZDGpD4sKKVMqrs4sjbIEwt1AP/rMQD2lsjBHu6j1aFdqGYxEe5qk1qQ59p6mWt+4pft0We2xyc
SpiaKh3h6OB2RffzeSFgA5mx29HnbMKod/nAgDsg+HfZmk3hPZpgodXTssKmthghHyTZX+4StCQl
jwx9b3eeE6uhNeGRYi6DVVYGhb7k5ZQ10F06l6PSPxcNkoG80xXihSwa39shL433Y7NfKBgjCmr0
NeGTnPvDo1pkAh0o/JFaJS3So0h5CGjqUJwoIOuPeOofwVfsmUmMloeZ/EpjMP+OjLhWW4nMCcST
tgyLuhJZ+HP/CaV74aom0bzUiWwrC3xgaO7zrSZuC/BxI/EKARk0k9T6Ym6jByVHyQ0QCz4z1CG1
BdGskSPndkxIp3Um6HJT0Q7amno2PfttV/cDmb4N8Rhq4Ytu68y363Y47COfPUw310hGKgBKpiOL
2gfgSqPPka2Be+V/9txSGhEgXhYWRpzK80dJYskUaKlQb7bidjdZqoL1zs4E+QIgxLSvINPlDDmZ
qxjGN7U8eyeDFY3U67T04VhvWYVZBkHNz5Yt9O/t/q5QpN9Zpl7jO397L2jbAK/G1ZmjEB4XH4p+
kj1OgWoGSSOxYh5CqDXF28CkjippLjPeXqZheanZIHjT1oVApnVpb4XvtGYFkM0xkQd0p7Zurc2o
7pS19C/nQ8OP6syUIQ617m2YqmuDEO9sECcQlxhbvaACJVr5BnetJfHubTWk+O0KjHGnTKnxFLPc
qiD+vYhV3Ir+fIFec9t1xvHgyyv33uKplGqLpiUGM60N4BN8IJQhKPH1UHSl3I4nlp8gjZ2idKi7
qMC7n9ffdnlBqvcYph4jpUP0YBXUnTpw7RZYQGsRKSKwlb9hjbTsUw0xltbdjEZog96UHvk3VDpR
CxIPgAX8A574LwgRGJLCJMMc4ob6Jyqp4lRExbqss7po3hQGiQgScr/2j2GDHEEe1VEWcKEbpR9I
Icfv7/O5S1N+xXtrZ3V+bQsrTm4FKG6wLhaeVVlN7sI8sGFzzHaC3ylS6VByDuSHLlQNlGfRbC83
fHkE5aJ0d+uxUSB8Bqu7kNSjCbpBMfGK0ZK5rert9fVfhDGn6qZMOhz1SvT8E233hyUM7mdIk2Sf
kwfD2hcKNv2XEzw2HdSU1aogy4oJB0vzgUuvqwuvK4usnlmXspcyYbRW98dMTDzlXeT3GC0VcLaM
PFEWspxiZW7QyTUylaP9kYIyO57IxyNnBw/aqLOxvJSsDiy2h97t1DLfnUWNTaSYQO+Nsag3bZLU
zuESR0NOjGpG9YYc2x2b6A/En3dmd/khHBYOwxi2jIYYmb3M+makjwrLSOy4pqzOUfszWfH7b9g6
qTb2UWC3wZBznGiJ+7wHOZo624mq/Bo1LMCn14+CtaoFaK8wkXQyKvaoU5gPiHK7kvewLy7+ljML
3UJPwinwaO7DrBbVt8vjhqhL9bobGy3FSWA3vcPj8dYE18fGM2lPh/JbxKc68zXsfiJ7E959bHW/
cUKpX6vCaJ8sHWnS7EMg3HpAYkgGDWY0QB1MaAmY0MUPQ+tK2FYhDYMaZtomZpXFOTQEVqO3AAgZ
C0wEQfGOY6c9h6Ri7D8ER5riO4XUu5YEJOaCxQw/5YHqiolCOLXKtSUkAyXmihZTJz7I3CGZautW
2pEDToQbc+HNy19Thdc0e9eCDusF4noE3Y8d54ruCVhAKkGF+XMeG03ZpEFBHA0zjSKBh6iRS++X
TMHTc5ICNXd8/qsSOiWYKj3qMB4T0k+WT4auFT6v5DIUdbJfi+sO5nP/jKS7DH7oCP4xf9bD7HVl
ECFWK68Z55X2AdvrXi0JaVusAxQOGUo1hcOLsydHrV/Md7BsMe7J17c5btb0K0zOYREIiisFTCHa
l1wXDUfWv2fHtIwqHzrUwJ9ieS1devLK38p4R+zec5xocfujcOXHkp9fC0ZOjH+KmH9Xo2RkHqhd
+W7QnBAFjG6eBCmwWeDRHq/qJh/wnYhTXiGybI3SweGG5t0nVOknXntxo3KgwuEor4inRXeM5yNa
LO4ajqUtf6KJpb+TL92oKAHYbSsYA1nLAlqfP0p+v7Hsi31psPaWj8DChrAWdtmqo6W6TNnwrg9Y
IgJGQcF4DEr8/07iTi/d1X2Aig7p+1n7vOiE77bu8N2ZpZ8VP06zybuowXVF+dNho3LJSD3R5M+m
86P9HiiG+FMnFnsyZ0SLwRxtC6kYygsz6ihVpWiVUSLw+MsRvyl8BNav4JiU6CfUEfiQKZtzwJih
F8LYBh1EuG23ylkoRjEGMxSOYWgLpqU3FLpGvJa+KZa9kipv/KuZM2BFrQbYHnaI5wiCt8PEpnKL
ZU1OwLx6ErttMcs8BWsP3bDsj72x2uOJHiVzYZfd/Q8jMQVKZspUUyKfJz1q+VoBmiYNO8AI9Wqg
Ig2QiTtfXvAek5PIK4v02/hR8On5ASaxF4ngLqHgIWPInKkn1EPjFOzsbPYJ9j6BXUbT7eU4i5JD
1IajpnhwdtsoUB16E6tl9HO8Bf6GR3SfiQAjZcKucor7GHn6Pu1ZmAQKCDGizxPCWcTYN4VFlOhZ
9bAJLnpGuK6g5BacRxYQ/yPeBDvYVuJSs2oMnDiPBFYHHbvG960tIK/IL7QQhCU3/wZM7DVMqSi4
Ih6aFOZKvqsnoVDTvgINwfIde0CRRtDBiZaj0M9SkAkl3xJkgWDH90kRGPI4eG/3tEBEeb+pChRS
Z/n8MQHvwz8N140dr/vOwrkFI1H10O9mj031219W9bMrQZdfuIqPu69m75d8K9aprwq1lryp2AK5
vpcwHEO5vAxrh6EY7FZNF4ulgXX4eJZXQNyBJ+t9V42l+o/oAwOudR5S+APRYBmOXFHawnU0cFpe
FJTHAKV562qtGPlmP8H+WDR18l4X/dBg34OI2tQPjGKjDD5QEeOK7gv1QxU2O3oeOdEX/H6X5voV
Q4qezxpK22qtPj0sLn7mNtfsoS1+JjsKNCZg9HKT/lGhgm6HhyxDchAjZn5TRHTHp1UZOO1ZlCPQ
5R8Oz/OO5oEh3WP0H3deVupNaT8+yfL2vv72ckN5IxJ/ysZwlTdvc8txN58rxaCBjWL7n3mCM5D8
d0pz5K3Twdx/JMFn+cFdV8NXTZLHVi3BecXcKZHRu+56IwZc8sZ4+s7OxfXX6QQ71RdOmkxhGudL
ypxTLlVWrVZFHJfVUWIjyqijfiHEcfSo4jptOpVuV5EkaTAqo3vt/maFGfdlwNJA2L1fJGsYyPvX
KNrwk/QPmyl6hmQ1Oh6u0TI4fIJNEfkbC6aipf7yf7atX/6b0+pL7NyNkpDsZKLa95GZhbqc1FF5
vs8E14CSJCLl0eBLOM1V6ywHOBwPzIlUczcnXiJcs7rzobN5HbGke7Sh/zd/mWgkUY4r1upeEZG1
VfvDWpjaAAtqmVwpPcw52FEKN53HTRfzS5IOj7aXIup5J3gW8onGfYUjQQqUsUgNeQvY1pfcc8ph
/PLOX0kyLKsUZ0d6RPPB+u36924ZY3HgEHPGjCmqkeNjcNmHb7XqdOMb++fK6NSR8WtEy7OEUbnZ
0my0cVRS/IK/60qTRSo86i4k51NS8PQv/hXrYYFhQ5/DO+ebpsOa1pn5qquMxqbmY+Yc6MwzTxXg
ceqbQCi50CcCkYkVJXxh7Rq+DTU7+UXLuE5bYk7+bhNz79JfesLiIKmUDwrq9S/RChavDS8Oide+
PP3ZlM+uMhXzoZay7rgYhhUBdK/QMWESuWu3HStoAvSkoP94MgQ/4mCHaUdKptNgNCSuFAueVE5M
dXGq+rl7VS+BaUjalAkcirhO+J4y7H1ycTaNiM5Wf188XvMEwgsiuA1jsplb/N7IU2dRIV0nar0R
6eiu8fgfKG3D2Ehn26RMl+ctqCAOVg1fM+WkGgexsa2aSGbwBPIF7mQrvxXTfPH0c3jg2V0XtjYi
Grd46HrzITmpfXqAQIdhy/ae8Wb5AF3ynXfmX5dMnd5gKzBRYK7N+CaxZAIuHV9eKDQOo/em1RAr
ItYpajevkbk6+gbtR5vLS2GX5ZaBAA+oDpDc2Vvd3mxvCqvmykD3F7L5A539zZettNXhewa6kL2E
y0gyLbHWCopWZX1xa5m7UPewipFrxttZljf32GcAPP/O5iIi0qJA5o7n95Kp62IUIKx9Kj9xtS2i
1/jXt8YDq6YoOEA9WNvcXAF/x/+/oY+RNLgCokAwWh9gVwdJ6wuohyCo/ruoHswccpkFYvy+IZuA
YgEQSAOhcjeuumhwhN5RPKwc8wighcuOuIcKE82iY2GCcIkpomI7I/VWW95Pu2hRlIW+QKUWTSvr
Jb5faGWwP8zZ3C0W7C/vVSavOPUd59lD7sFHOilCx4fBpAXSR/DK1v05lFU3PZw1YTfCm2l1zDQ7
GThYJdg/xn/3ov/OwBP5xiVFVnuHkhitwseXjX6YfW01pgq1vPkhCmT7hOrGsCjbWyHAA8jov6X7
G3pGlp2LF1AR8I0UCD30sjpguahGI/QcYCNDCwNK3TglTDvnuSkmyJHmB/6YLTMsseKlO/+R8wDp
xt57s/kkPJ9llENXGKjEuWuNFZJGXtKGsOFgyjTsefTb89tfY02xYJX67RiK87MPso4N3tCszreb
zkg4b49w7GOYBP+epexvdIl+kxtcfCPY2xQfkxvAZSC7VJW9GELvig8CHy0/Zlq5BbUfslkg7JtE
2pg1WWNodDiNDOSTim27bckI7LKU1OMT4rirPGb+xupmO2FHZWAR6HDAt5/2d2JPozsXRjLjukUm
GYfguT8EjBphsHK4gwPbjryhwDGw7MGSOToE11lRLB4SH5l4X7MycG5ryffL54Fkm9dZRLOIaXGX
I+0Ah/O3OUIoACZ0Jtp6qn+Zmt9vlp3DvWtRUiLKyQQsevraydH4a+tRbWeJSO4gbnoa12bezwBU
hjjJLHF7Nht4tQF8FsEuUlph6EDAj37D9IyhkDAoLSTIaCBSZdsrWroP0UiX61krS4J87zmmw7Mp
T1Rc+CtnF80pGFwwuqOOqgrxSrqkq0lYCb7U7em/CGG4PPWNw0Gohdo4TpYOD0KVUfyWFaaigStW
R6hOGcAvGQQYc2AiLilCMU7wbEBu3TyyFYR0AA60bslbzzfDY8rDEM3sWvGbLQSrJOeo9MabWqIg
wEb+bzZQ7omZkbRUaEXEtqvFN6ofDda5nkADpveusrDPpEyfCSuNdv0QkgC52LaVdfGi35r59g6I
kEgPBB2J5LN/ow4DAB2blcI4M53eNBKAcmN6RB8SRqDANl18SnwvOcgky+n32/edFXF2YBHPWqOL
v8WE48ejixVDkdos3GZeq8X3JwrbupiZLJbqb6MJwJ7YvMJRGCWoCLrNe/D2dNZhQ1Jo5gCJSOeO
CTIeS3VGpLYt/JtM1TG6Rkreg/CT8JoDaJcfGUaToS2nTIoDBQ+jcHSr0k/7Qe6IMsG4ZWOKT4Qp
YjIW45IFIcYBJnpXlegZC3JMDQHoJ/pT1tersmp48Yu8v0jA7BKBJqXQ9OvxV7crvaFbGQExLcMc
RlhvijaEuq1AHDCVGy5ZyfPuOm40bJJZZqeF7aHrhPrxr/KQr+sldV5lzubgqQtb1BoHAANp4KpD
DGpkpTcDO1yEXlPzbBOs1Eay2M1STv85sOpgIS7FRiF82Mmt5WtGJ+0MNcVAW4gb3wsSHRvLvIUX
AOcQMUhhOcwA8IyEqJFxoGsoGVAXwj8WI0CcbFT5KTSRrD2TJKIsWEoZ6xWpT8zOWVOShpeQ/Awx
Qi1n4B/zhqNK2q8E73YBMDyotvFno8WP4bE7fInPuXtrRAcBeTNsWy32JXdIFu+QB16CHVGMEHEM
cVQSNbgiHB28i7KjmDGhTq+Oli3J1lA6OzM0Ml/wKDwX2MjMEyRyu8X3qfAV4I2n32Co1uZCHJWt
aw2etiuSks3MM5soCpjKYuLzYpOYmg3JMPZdyKXKiaKvnOKs/R8HF4zXCXgxdrV9EkuO5tBDHND+
nmZZCtEkV7zSVy/cbk+Sn/ymfvLqhcy6RYfxCyDQESH1VE5+hNg8NgGSLt9aJGONF06qMOKaoVyw
QhYY/NZJLUmmc/Veg9xdKab8OOuG8Bd/xqpPoxLipahmyw0m68IGg9JFw/C9K1IKzPedquYVR/pC
mB1+yWXFyJVSyZN60saSZG7Sl0ZyhpZBhPIIprugdQtXV5I2WIxkgnDWXE2t3cSWOw5IB8JAGnqq
MkjVahYdOw/PIZmtlxFM0nfj38QKslyKFRE/oJPImujOBG5XPTSnKKHPgNItVex4DoD6CL8Oc0Ew
dbcQ2GYZxEFl/SzYvi+0Zk/l7MIJpVF4sgjyjPniHoJYNSBc7cquDMLP/OR/2KyObBBOrVYJeGD/
d7YAx3kpAztS0pHr9ol7bVQHSsdPPfnPWehfUSosJTEAflMmkRAPL6tasfucvMmaRDX9/SxqlUJC
Pmxk1/SCcHEfVFwlpTN48nzJ/abpVxkE1gJWYSZllcxgnhT6zvpKEXzAF/1/mT71bUeX9CGNFNMf
sz0I8xvjnDBRcK5GM5HMq3tcDbK2EDCJrSXSX/KEyKK8d7OMgL3XtU5OYJTCsj8+8zn1wYvOuk0F
sn3Qxa/aMAvGPQ0iLW3k+ctepMjLnVMgsVJJpYVHBRs/B1sEhwoyd9a98cMLusZ5DOz7Ooqd+PdK
Cwtnt9nWbdDmvjlBTJATcsi1FT3Z0JEbPMQoSvmZKaJbkGZhLeV6iEe+7g6EJJ+1bg+QelWkrPgx
Xsu+SZLx3KTlE/zbfRIsD670EdpMDv+J6cjmVApOXHdDHfM+xkJYl89NvUGdSrbbSpnk/Kbe+dbX
Lj5mbY09txhZ2d4aRb7zyXBsO8hoI3qUBEx4/JwA7WfcicQoUKQOL0udHHIM5eqlskHRtZEUfOp6
VdEzQuP70WpCT63mLvmASVF+M+IpnWGZYgkFek1a1Wi/VKwF9ifyIz/ZqZQJUfcDe/kp6ZWcINhW
KS6EIKpJcg4GAvMJTe4q81o9d5VLOWvKpr7jhogYcsQhBZKXeAn2BvU1TJ39MjoEMuEXyO2x266x
DGhnPwiXIVKAmjUOsylntgSf+PCaokQAPqi0n0J0crp7yLZ9mde/uGkmRY8D52vu0voOWTYnEzBe
lspZGokozXKYTKdrld1FVxIk67t2uQzQRtMFKGU5g3Z8dmQLlXIz8dIKrS2gyhPniYwBQWbahRZW
UzgG6GJloqyamlKpmLRIS0EO4SDMlWsiE42Ig9Tbo9ptGKMdCSxkrzXtUVfsB4XWQJL50ia9Kn1C
AqfFvQRJaZk4WBSYcf5IZBjchzxrHHU6E/8LqKGJdRk8lBAZ/8gyd4aSBrCuqM/78aMYDWldo7r/
cI42S9Xb12tRvByvNGBfFm03MYptolTAh1nAc6jLPO96qgItH5KfY4+r0nwB51Ym3lw8pa3v61U2
ddSnZOmcFRSVlX+ZrSpah7vF7pXYweXg5681qB7VScjwqrFpGMRCAezXcXeq4pri4YTSTGFI65aQ
g2HSqXL+jXg0mrx0v5F3WGx/NM8gEzCKrjge4Cl7hflLM13pKCzofUStNok6vEJVQc9lkJWMXYJk
aAb+/kc3SlG4ANBmpk0vxFjlv9fA9et1s2qLz1ERyjkGh6zqMM9tYCVKTOlXkih/Av8wYk47bcla
jGCEUI61quZiwEO98bOx9pmgoLEZqU//X61K5MTLPm1p+r9QERyPuJ/TIW0XppE1dY9MawEuOYFu
wglkrgqqSaqpmnsuJ50+2qgC7kxan/j8r5/0icimBb1pIYKG8drgDeTE6Ssq6QA0WC4e8os9nLjC
IcYReS99956YAYoKULCqr8LTgZry8XFHfso4rHtOfLg4CaEsONqzs4T7Y8qPuefkVzM7K2vyJkzQ
3URw8YW4dEuXyXnRLWLvjA20YaToSlBUaBIvkSCdttVm6kAHar4FQD/ZudpBFGPeec0t7ZlPryYU
jdg9XDucBgDA2gFXYt4i9FZEXrNdkvISS1eXNQNxZKuH63dD2cT8S/HQK5jJvIruB/c6ehyJsl0y
nW3SjoB+GVp0YFRyOapFTNDddgpMa0PcvmfwIfAEjM5+1S2Lm8HWBdmFDPEOTBdTgbVuC9scbkPE
wy9BhnSg5LNvD9qtWcFRAZdgb0VJedl8EyFUPMobZ/Ag+ncNlotbLb8XFLFjAsc2tUk+q2KOUF97
o3wXl05kj7YxzykZGhOVNRqlUnXzHE83NmwM4N/DYF5EOB1UpR1ZKmw3/d6ylCuhiLDP7aP4Tq9R
96gY5vTUrEGkF08bBnW0rhbpOPZ3KqqDDULB4Hvljg5tP0H3V5SnW/sp4Kly2VfnO2jTlHsQiQVQ
4ERqpmyOktlUJQ0w5vbztGJsvsvxcYcE8rrFYIY9Oy05hbF5PbjUQ0jIeIi/XkJ3CF9FXk+S+rNi
IPVrn4v5F3KS3oz4knr/YMk6Wg/UVhAxyxibPm5fuUGx9zbgFw43TNFf7bHMM4/b2EPmUoydXw3m
lcSB+jbi2P7N2TFbxGUqzD6nJ9wU2FtWfSPcOwDNHnVMJnTeuJXP2eUaS6zR+Xxe3PAWeSy4HPhf
72y4yzWPfUuWTHpWisQ0lbLl7Pj8DITr7pKG8PWc+/jlUd855WXLKAYjvX03HoDi9XV82I2a9umw
nURCLyuaqtFIlCYkOJ2ZY8jCuRzktp0sLt4Xl3acIc35FYHsQVHL7/5SITZHozYvXRBVxtRXNTen
+bRNwD5RZr5dQfWCnYhApSYklRHwP//jQCrL5MleAXgMpupRto0rXHyTicX1Bh9PM4tMzxYsW5rj
aKpKML4BfZ7OJDCxmC+0u1n/BxXXMBjfueFf0cxjr0PTmXfRsYOiXNNnpJsvVNJqVS1x3JdGx+wp
HLwrjP56KAowqdTXJL8ObskL8X73QYPh4OQWftHmWZIFi+E0BDmhdtiWIyBzFn5h5LiantCyhE7n
49bdYr9aYm5Ir7VPSue2+1/yc3VMDtTVlijFLml7WqIyI+dnpAejvpe3jgsyj6BnwzssJtPEeul4
/ODIodVqkpqG7ykkEhbu9LBW0ZalmYT3Uyxm1C/rBSLQe0eoAgT9cGeyBvVOybewMnVUSMoqjauJ
Mg4U0SMtw2y93ucFDs7bj/X2dF94rdy6ZcEk/vDaf7aCq5DA2N9Un2fSEfm6mzNu38c4GDKJnSMJ
gC6+iJSS6ERQfyTLpxEfycSMMHmAttaqFi++nT//M43tUceIAXU+AMNzAWyNbKBfDfIDa8+0MQYP
x3ARMP8whMq93j/cTiOMKCSN2DsvaQfP60LAIYhuL6HSSqqaMEvQ8Wmm0LzDnjAcF8qf6k8dLNVk
x4mHB+rEzJW6XQ66i7i/Itlk2RgDtxWTcQWU8Op/oNZUzdf3myjaWLbGAIc3uevVQI6t8R5UgfbJ
xrN08S4A+6jdOGAPHMsF9Z4K+aYmbZU2Ng2OmiXHNfZFUSPdRnM0f9BmvM7qxis85xNlfEJEHAPL
n0Zcvy/TmA826y/ElFCgi9NmkXIFE9I15TFvjqkWZXQ9U32Xo/lhPQOK/v/6TClFhvLieiNqapbS
XJs9tdNH4vJEEcBSGNGuaO13SwYoWiCwGKzd4V3Yt3R0cinXk5nlE0/+lYTP1tc4dEbBzWHYZ32p
RKuF0GzF8h047bo9b3cnPHwaN+/Oyye8gblzppgIIl/rKwVIrirg7hiSu4W4YBs9Jue/JauRtT8y
vUA1OgL0z/C6XsbOOw7+n3IwgIwzjmfYDQ9BsB4y5M3ckz/ErkrsvkQ6zZT7tuzqBSj9kUaV2Xi+
zLpzUtFbGsR/w7aiz8yOYvcEqBiU7TLfIRF3Uv7ifjPKD4xD2X+f/bu5zSni4oXt5irjdugKcTjA
GDGacl5tDAvG0OCueXToP1at2CLhsK0dv3cHiQ5Dv9aZWHceJ8y5yYiaTvF0LoF9UNjX16EMcPcm
3qlLS8t03G2GXBKF2tv5DyhB7nUOqOXsiwVZ2MkTZMRXbbjo6woUShCJNVJylFI9X2D+3IgAA283
0r6GgzT195j06uZFkyfnLkn9mWBgJDzyhh36JvWXMyplrzcymoQDPntE4iFTX/LlSb9rf4FY18Tv
771uqw0t8l8lglrqN8JzabDxEJORi3AyvwP8HV8dIKyaRrO+j1ixO0gfR3IHAGA0l/AlzeFSUqVH
iyfWpy2vb2MuecHUuquNCqq/XcchRP1Oc535jVWMJhD63VFfY/IQ2xbevtmm4AZj5JCeYWv/eYwt
jmAgMhiW1G1bi+c0M1W9qAkK5l5vKiUQ44JuacKF0hRNGbwMwVHb9kmrbVqPiqs4qsuP0YtZqpNw
wNv39FPWcdtOS4HCy7aekCqo9cntuKp0NU/9NjD7peRK1aKl1rqjPSvh/8swL6npCk0Try7gx8kR
LTR7gCJbc6/vE74k8j9ePUqtVuLexTbAn5gntfbDGwjfO8pV2WuRkdAnUytyVNGcsiHK9IgjphcR
qyj/ILOMDhopYs4jnLRVhcJU/jZC1+8bF6hGhOuoeK+VUe2lG5A008ThwAvHGVv+nhbL+7YD9VJF
cgM45+kMHncdz1tyzHBkUI9DCNN7NdsskC+hbgIPf3iltcLXQjffdwJBfAUjQmRp377I2jCM+kdV
om+qjiEOOLnqkb1RZ2sW7J9tkU8RwCdrMygW4WfqxaedHPeK9jgd+dqylIMXt2SiKuxBCWQfVGh+
LwfkcDI6gDBRdF7o01TnKwMY9W6AxYOgjy4+RKlSMlyqPom4VgDqyRzmnYymJitTIlcQYenugKBm
I1p4Nr17XVOEYsbusugCwKu3hYM26hCA4c7N6eLRsAZkW4sDXA6MZbAH2kflNpNkg2Z+7czBqjjd
GH3a/LC6+zNxrxlTYQZvRpHpa+bfZulOxeshBfjMBpkRBZ/3M9Lrj8OvepZfQ1j1XYsM/iaJoL7r
KhnMtl4ostMIJKKeFR44uhZkSRwtoJHejkJk2Q25kNc4NO6j0/PsjX5tgkR3OgCYl8IEWZ8JSM5G
37upgAFlMVsZlFhS2CWgs8lnuaLD+Zs2+yD6DCvZCoWIisIft/KIxwJZi4fuBEkx2jsqg2w4Vhjd
zU/vpxBsUFSEIwOWBnz2B9nk5E+1OXM5ygfsgRH6qBYg9FNhlPNlJ/EgGfCYxfBzDX1NYeyq+Ksz
fP3iR90otQi6sl2WGFugsQ1zvhjLiAqPAh7h+e9M3XDAOFbb/sy7TyrA+97khH5y7GDn5XLwbbFh
FXCPQ2hotZXr8E32lQQzUItImpu8bNbjPnoK7KqNqDHk4To3Sr7iVxUGBPmT8FRYgLYlTXran66g
4hNDeJs2fHgXUhXDE3bLUJi3YC5qopgvtCPMjAarc73/5aiVki/vcb50qoA/7IIAoWByMapXz4IO
5yPZ4JaSWk8Fq0oIru9N6L5LtEh3AR21F5i3ljOGh8Wz6inWVu+LFQ9jKGEj7hlVKP5cLFKRTOOM
fR/TmrQJCt6qt6QHiKnKimUm/6mbPRK40RvsE8rNkVO9jgZAejOs+QfhrVy9cw5aGHmSJTRg+yaA
9yJcnMnaXhY4cK56VJajlN658lSPR10t9dPxXW3w8dF5ZsowedzZ6S8STxGPL95V/rBDt+Iim0I/
I+1AYWL+YXqYTmbBUV+QsG5SU7IPXK+l7jTQONqrWMzjK0i0mGkmvRcwrG1x3cGKTHavY0PPYDNg
4F+oPm5LsAohAwdZr50WHmdnr2WpBzMBCRXKulVtO1pU8MKxCjJC/i+l3CJ03x1QY53+W3UZ/d91
R/Hvpe25l/146aZDL56RJ/+omSHSQo8Skg7MSBN87IiSbqGKY4grLzKJtyvkuc/n1gjRFH+9w7Hl
7yvfxQv+d9Uk9MTocWsaz/8xMkehbOi7dYTF603R+DB222373XrwhIeKCN51ahGdANEwbiVW8oTM
+G78Nm/Mdwv+xVUjJkqHQPPf5ERYtZs2wsEnjIMX3jgcFExim8JmeS72OKcHJ5b+ZO2kq3X9sNBX
T8d+H+pTXLLBAJ/jf4qr+UItxRNmL5+Lp6llT5R9AybLQKBAOmVcpZbLIh5ND/90vtP/NXw5ncWi
xr9icOo17FVFEC3GAWrYM/G/JCYMazObsAX4lhr8pFRkXrfxv37hO5yQaD6bo8EcugagIODTHle5
eqIeI10XEf7L2fPfsufeVmU++Wu7fs54NUBRw8g/rReNx7zl7mCqacn3H9rXNXzNUi4K5epq9SQB
IdLGdGWPlEGVHDC0BiH2bmkoKFuFTbJJwA4Bw2/v6X+oEhCbGRX1Ny3a++1DWDhM1y2UXmppvMLo
ZLCKilxozuxrZ0EftoMFcH7yYhTxH9SbQ6ngbPtptu7ARp5tcPBUWwKJmfWsSDxCqhM6VJqepJNx
MOVYRKbnduGI6nVd409PyLeiexRGd4rijsU3MVMXWE3ZOx9fOmH6dXQPH/vahy4pf7I4LsfV9cI9
eGta9BEVKUJHi0vt45RtfWElE+vkC9IXPKOQLylCK2KGQ/Fbs6DuRQcJavq+8GwgWEwF6Fi6wauG
0hKedunhffz93SLrBmSIDXFEis0D9xbidxzEfDYN45iBt/ET8jdkrU1zKQRmrVRI+vQqK9xrDNjL
g3H/d9Ukvif+SEIfCZ/g3WoqEz7mlHyeyfOpenbBAAK2ivjLZfLWRZo8pw5+8hc9SEUIiyUGeye2
O1x8FTBGF/IGktBS4HrOlQjZ3b0nMkyNm84rwGiScqBNyi7hiwQlrGLLAm1eY4PTTIByit8xWatc
kOEQfkXLfNt4mkwwe9Rp+MuOLzLloPieCLodb/wS4/AidNKZQd/dbFAHx5nHUAOVx0GbtyGGO1jT
fm/YAUuDcjVrF8T7O7FlAqUo+ll7fWUIjltyyhfj5+bpd0PRDLuLro53mwQT56ss1HXwX1C8doWD
euUxHOlXwKpKzTp5UB1hTWle4tyG8KjP9zQA4VMUHrNoOHkwcD5t4adCmNU3bEM6SpyqiY9SATO6
DFjZk+H1rzmOO823ihPq8+YN0/MG+eFqZ5npzlS3V5N6hLEk3dGGxza1k1hvbBB7jI/ZFMK5k7RG
o+ZtDiU29WB8uvKkXL8hihCYrH7VSEFL9KIrBRW2kaxisIrNRK/aGv9v0p9QUxG6lSvYEAZ1oyax
X+j9aTYuIGYXLBmKVCiaUbGxPiEKivd+M8Pr8A/OD/6caraf1GIuLkGg+V96wBjAF4KtV2D5LB5d
mIngVSH1Z8jpl9+yz7y91wGr1c8E4hrUTprsqWdeAdoDuwNXuT/nsdL89RzbrhtvDISYPtdw8G7N
DftvVURbwCKEtdQHGbe5x+XAudXDF6vM2u2wzNXf8V4U81UYmkOxJEWQrqjcPMtEAPMJC6VITWAo
EJ8xVA60BOMxkJyWt8uokj9EIEA2nR1RQQDY43Ezo2DUX6Y1dAjbbg1vppgP1mg/vEqESfvRio/5
g9su3j4huWeWit9LR3LfcYaeJq4dxMPdcX6NICJnYGetbB+WuFKpbqwupm7PvOaLtndzjf9LSmjp
G3sOilzWmiTmZr5VdhTKQh2P/u9MUXIfnVT2duOlWHhSAx0Oe/VRUZWWrB07xcGiwXa+o5q2FpFD
bELBiA2GEZpGeyQcB4TMqPGMQZEa06DhWoxQEvGaeei9B8ZieFrFqlnfDVww2Y9DRDoeBdCHGFiD
yQVSrFcqHleP3rh+e82lXwhVScc8hP6PPUC+unF71FEwoodLQE6sBNC9pKEC/TSbPlFjASPz4cq5
tGEdPD0sT3VHl7Cux/qlR8Yv+sBAmCIwH78gtMgCRQkAW4gQwgsSHDlhNJF4ipVqxi6FC/EegoXd
udIlmPsGS7onRIWGQkzynIvG8hX5/b2SpMGf26IW4b52kuGxg/cbSG4etwtQLYmyvn7gMimx5Tgt
aEoAFEFMs7Fz0J8/9mXgfBbV1wzsHF3XbmR1A6NQa6UVfD8fsp1LU8W4LSXjc2BXC/1QnwA1ZEsz
Kr117qHQrOFBiH93Yv+FyEmxP4irHevs7j7Cov+3uf92tXgaZQa4NCn9C7XhWLeaqpOoilM1fgCE
3XKpwajEmbOVc+EsqalidRbpG8i8C+Uh+eth7WtJdZnI4j0zlc/m2P2cgdBwXYLa3D5NAAIMj8SR
mZkkTT/Uq+kvOAEhQQDdEmljDk1XGAHg55SnSFPIt6ILx75npizHLEwvtH5gEhtuP3PpcGE2bZv3
xgQSwcbvdzQZ2u/NIZgcatR9zelJ/rzzNb/lQyPn4Zrm/9/F3PRGaRFkvuC8GXmgu6bkQppbh5pg
IgM8AYuO0236igJubylTu2LTw9yYR7Il2/p+540edK/n9+di9amOd0YzJ8d/24QlQyLfwyRtNG2f
tJGW+jFoSNfhAXxEyGn2yn/Fn7tMlkLZE8FhoWaEOuaRTevtxtda7mNnIQuSuZxhppM2N8gFw04C
5LOl3nuEhzyPIq8WuoxUNHKdhdsfXsDlrG8lI3MtwEiokxSZ6tH+l+aChU0ZJa1Aw6In7EyBZKmc
Jgvozj/YMzGkraTtesPMAucARuAfcyTl6hBMBQmmOzlmehZ1hQfKQBymi9jRu9KwLqYbSY9OY/U+
kEvtSe3cIa++QzfYQgl5L8KMd4IxyONc+3RGA6FU6/LrtePLB1Zw+2oO/oyVqvbbrY2IFoJti4kp
s6e2igJ+0ntYgZbnnw8ukI91Bn0gr4KGhjP2pLoMA4jkYs1MgmBtpFxhYgaXY0EtbTr0vK5QVEVt
fsXsiCHRnJeT97XlDnt5OG0+WH1SbowYAGElV2OJukpT10t9Tuhv7BIZf5JT5QWc39nJJANqTLvv
MxtcAW4TAgStnWWzmrLUabEgrfReMV7Lk7O7fYP8C6dHoQVHviP66izOCwoAZgzj5uTlGm98El8z
7IEvE83F2l9lmVlCXxTCly7VzsND8SEmvpb+bOaAvZitjIfXfcgsIyqKo0X07wL1WC79+bNo0Io2
VkQaTG6vRPqD5QxOWs0+YbPSb60dT9ANbnUYQQAhM3DPhg7u39vMx1OUuYmr+g9RjNYodSsQlo3+
pZpGzdBDJOeubB5IizHkUOFD6Fp7BDkwA5Q7IPDZJeFIiFgTNRZIZ9GdhnqOecOsuUNnt5Ld2bUa
lnfMMhKdszR5CWePV92URCE+DXGsCvILq7oVubKUnjwAXf8r7Jx2lbUeNGNesygYSIqtqd6FBSXV
Ofuc7KgT2HFvD3FS8ouUVsv5J+/Mc9xxlx1lr3lPIVwd3tfBAV40V5qofM6+eOTJ9XiUt5XCKX/o
i+FjXaeZ9/HcWD7GQmDADpqrIS/brCuYQKyyqmfb/PxpeNlb6GB8x5sL4WvtiiDHaFT4Ah51WmzM
cweYmmS7b9N7DK4VRuBDmNyelilOlfV4uuHpjQkmwtuuqJx0+ZZDVqP4DoSYRT+t40Ggqpa47aOx
y+kTCoEB2lIgG87FkQK+mGLNJJTjupMRciQjHnJNQEqO9uFaYZE5J1bzQvNZKaJPhyD9D4QBCsf0
IdRc4oKa5MFwVeby3b0EQC+xsAN3catmSQeHuJ0rQZEE3+Uj4QfL9vhGbQD25T4C9Qc7fYTGWf3w
Ji1KkI8T/3smk1QmISjWAznBvLgkASzyaNTDF9w3Ye4LionJTgDbiBZW4+pFfDzZHtaWVMAh1IXR
AUE521ZhJZuwXRAFv/PDr0vAd3JzVrJtT8a254UPbnbWS1SWgLZEFD0t7Xo/hBMS/DY5GAV9UnSt
1ObFowmZ8eia9/Q883E597o2NJWW2p53NbYRyY3+eeXXw0Sjy7FSmS+B3ZE/y8w6Y7gsTIlEE1Zp
oCrTG55WvcykGof8xJmGlRdCmIkuVy5xWpyG2Wgs4sr7Ii5j4qYedH4lfCdfAJq/4HIIz69tIDOQ
yIayuzFes7IlAsfP9D83eoHDWcKzhpHoswJyAZ6l3SYnt0fjCXyVgqIFfaiDxGRmyQzLDGdbydWj
OXBb1NcloUMqPxcfVXsrIfhLiMtFbJcIDqZCjdflu1ADPCtYfPgHEo26TZOBL/3Qrqc2wE8yaLJs
VBsNEofMlUI/tE/c1nwfYza009hd361fKgOqziBuvSAdTCQv6jN0+ofVL/4QgKPzznBmPN6eqy9k
DuRuBUsHgyJP6N5a9HqRaRd1mmhbEZ/G2hZL8OlYolRRY1vqODDCbLYeSUxXYSJ2vbQQ1nhz7Zq1
yPhXo69Jvk4/sdD7ZizDDA7gRUyan4e2vTEzdeF5zrBCEb6n7a4EnOA7pwb6iEG3EDt2JlKn3j9N
CrduJ0A8etVMQHc1vpBx1envmEyQBuAc51mb2mXCQBsYtjK783gK7+k0kiceYpin4SfYxcxMhDNH
i2OxtFBk0Hi+kmvbiQGguccy9glZ+rOp9w9QeBV3Rd8/x3wFJRxdyDOqydlVyHxXeE53k3cEhRFT
gu7uUC/b98SOvni3ah51AFasZMCJhS/gqafRpEdSpfae/2e6D3y6OvwqG9Vt5H3fWULQWqYh/aI4
mGiKrzbW9nTFXc75L+SKgFF/iVyegUk97aokKMb+DfyF03+dy3Gr6zOpMncl5C9xefVznlsQrsNi
7uJYJvwfGQbYxC92IIZYG759TvZ2Bxtt+paToSoiZU26p2d98NYPTjtQLAcpvrfkHD1KzuFG/OEd
JDCuaWPfN5zW2I7ji3fYhLeHC49z024aZScoEEcBX6fhLgI6ycBpBaiuOFC0hVCdgZtm48VQyAXd
gXgsnPBpJYn5fRgtLZJxey145XUOjcxvVbAamIWfBy5P3LW8HgQN+5kAx78Nd4Apn3e71aN/kCft
E5GaiiAr3sWZkqSaZb7LBQiXrbrcv8MzigYFg3Thb7xJx3/nBb46N7Pv6r5IxpQwGlJiNpuVk129
X8UubGuG7ysMCixSzJf2Ol8ZdS8k4zTiOwOSvr3dsUVxGFnZ8Rh/PHRSKGeBe8sjyMqxwbZfwam6
rk3EPuxspRbR0kj8q48no1SCpuDzTH4jt3VvRLs26D42zctcuTzTbiG8YSXLkn9FY1X6FoXc5oBG
nBkf6WXDzufSAxnnSLzRmD/AMYw3GblDXqEG7XQmstERNcOGXpfT9cAQl13TUcIP7g0G7N26jozt
GDsPrG7RL4OCGIAYZ/zr+UMtyeezk6d3532PxLVYUurnSfopwsuBFSJ0qBZEdxEv9JeYEjT5XNZ1
L4YNYDvnXKPMyp6raebHkK852CAXSrQjLEDz8pUU1Gz0e6ddGhzaPlbHtaOc1o0UegMibONgl2GT
jMRWTFfDHkhPG32lGDf5ZIpaOyGjcZ1GiBm8jyLZmZVQWia5skAV3TWmuq+2t06qT0XyTVCnf+I9
tKiwNyBCfMTVYOifwWIBlxvaGy0YbaV7iKvBhTsXy/6vs76eHV5g62l5c9ZHI4qK2R2e/px8O1e8
d+hCqY8255lgYfoQpIgdGG3ijGQ4Dis962khp6MIMYKiovmqNZBwvClwjv3RK4XTyiKFdlWDYllJ
UOPxv63w/S1Et8R/4aH0afrGJIR/wvAv0JuhrqeS9GqbtdD8dme5/v9cNPMMpsqKLlRpUfd5+5qH
nsxVj+Kmz2+YdIsU+6iSlZuFeIvtaEHub3k2m5MKNypek84Ei8dyecc9F2TMVME9khRltm0y/1uO
dse8/5Qr/nYjU/wuSXvj29K1ej0lhc9o6ZUJbNXLifD5RcqPqAk78ZsfgIMiGEuAvk3795kggucw
noNONkySvLimL6tTusn6SWdoVL30WnjZVuGbDHXMK/IQDvdAZdWNr9FjzEy5Zs6vezLLCgyCCSxJ
JT/QTuagsLuxelLMB0B0wI1VWNbQARcIjlJfZ4izN/EEdwGs/xSL4YNybtpa14qcvu5EfN3z5BWt
44bMrQwJ27dyq/RV3goLHekgKpJoMS30M4boanziB84tKcEbSXT+T3FXYt4C7lhly/0rasXGVqA/
2LGgzeA+/VSvqQjSvBUAuORZQIvohok0O+dvzFa5wf1PBhqtBisAc5V94vZiGlzs020YfGRXRj5p
xe3cmE4SiAq1Yvv4afLWfc0Q4WJnOYzPZL8R/k30TKfYoXid3cAZ+lu2Wr+odEidiSXF2m2EvNKk
1xnjAaSa90eDwuNFNXP5Y8+OyDqQ30CoQWGFcHCX0c2oC/Y7CAvexar3glsRDwa7GWAc0Reb97Lo
DeatGp9mkzlX07q+ggFQKt5bNfRzIydf40+dVOEmv2CzCBpjUcM1N07T0oM6AkgwzXU+PjoBZsbj
kAnSd3pXbuYYtrbQKlVM1AG9CL/zpKifjCvQuok/MQ7PAe6uny7MDTlotkpxPzS3GS0UrJ0PzRPo
06iRUI+l/7yMNKHIleVqXKuMYkT8ATYt6TK/xC29vWY+0DvTeZKePj8xQ61WIj4Fa2ItsbOBP9Ny
BcwNysXCKDVzNaipMOBX6eIC4nR2Fpq4uXDge3Xf6yjgsHd504g1xc/AxPioSeUXjaVSWmMEy5ou
UGWb+3Y3CBec825WGHdeZasnte2mM9ym4yrmri+qH7Aervbypn01ycx/5G2bl/c+WlLvy54WmciQ
LGSwpu8OZ5l6y0ylfzcdHLzqzTRgtUCtvVnPDg5r8Zq2iYxt+4JsWPj1SDuv/0e0YLpVYJQusLFO
ckPxRk0fHIxHVO9vJSzGQBy3aAPXKFcI6PL/GtRZJjC4XND7NyLVof7CBBG0TF2goybFY/AVKzg9
ODOw+qzf0Rgv9Un7gX/c9+2d6cJT/BwdLP6ZZ0bCOAb62r6HIrbVDVjn2UqAkm4tr6ndGUrufALz
W+5n814Qjo42LBedpZrvn9g/gDZpyp+IIaiE3Bavf38L/+bOSmmTAdPHIIi+SGKoYnMwUWrCnB//
bYcoZwlpNy7VpbUoWQvGUkPFpsQ4xapa45m5HDAYlDfCBYogAdrA7WdzN8aDiS7gDw9dAZvMns5e
x9HrDRPON3r0vSVjiJQjRVJd/qIP4Qh7ovemcMT7EyhBvO28lzFN7fKuZMfIxQwYjNYAMcxcKr/S
cGFjeur0ZFPCS5+lMShEkeJl3NXpLW0LX2JtOk1EGMhU/wf/C9GLggrhrK7GbQY1phlNB5oHYp82
0hJBTYh1g9PoDgbJihgQtXudSua6zOleUxUkFgqKORP3P2u3Vzy37m5bQH2l1xRRJCRrbd/XIgSU
N9AKihnv+p+VvpdScmQ69pwEgwvwTdCa69uZ/lJKywM5RNJO8mHVeFK4GvnzwhbD0/0QruQEnIrY
Rgj7elfPCe1iilL3NFWwyr3tAgl0e8FiP+nnCVv6/mIsEX00tpJrQJmfcYrqMQvaBqYtCZ2XPts9
/G6GS56pGy0ws2VMD98LQwwW6SImHD+9Ya/q7zO2WFt+sWa7/fg+4m1ZQYpudwEIQHwCSTvfN/Ut
wJE99lJrPrADkDkE0OCy0tqXR9Q1J4MFQsWrKZbWc8v/l9439ysPPlmmVh96x1G8dqWAypoc3cPz
uH+J0DdjqRx1Q3uja68PQAhsReTmghnnkQgL/FUmkvNpX9NeDBY7+qQKQeJkHLCumPg5gW25BlzW
CReRPQDJR2ER/FMect9++N7aW1eeDOWxrMaSfBPZs4wqM3BATEw2Gms9fRKtUP0XqKOkGK31CVv6
u2DLGvQTPZISwYUVkxGd6Nqj8Th2cssgs3Rq65yq9xxr1pnSMWAefCVCAs2JEkg7QtOR84pFnATL
TJpumbieGqYguqEWywh5ITRJzCYUgW/NFYDIRyuu3K0Ix/FI/IkxrhXEQv4+5NEeLSWmfUX1BNpS
bb5YUeGpiluj+xZu4/zbociIPJmIcOKULEflVIsx4JamfIF6XYTZ0c5FmcgmTNQNhjM5yPmLpc+f
fGLBXJ1OZItZoZBog2F4wVhUKgeh+bOY0sPGZJlKRbW5uj3IxIYjVrRD+u8SFB8hRWdZnIM+RACm
jy9UvPW/qBmMXsu4oRbzLzFDjRHF+NtKPypqvT8b4IJXoDPwtgn6f8K0wKjTh8nWYfKS5tmEMp4S
cCzrW0hFkhmwAQJjEpVtdFX56YfjL5zhe3iGcT/9Vu7UgNkhX0zuGI8CIlmD/umBXqeVMMMCsQ79
uX+V5eM4n5r8ZRGNgkfVlMwu+pW8zr+8rD86A6LTvrCliF2Z9hgL6E8wMvLI4vZgtZBsfjtP+fbm
oDIKYT0/ZT35xGqsResTj8RsSPTqduTgl94mIh5l0Dohdw61ziWYb3dnLwBCWLWGrOvjCn3SXkv5
U6Eb4FZGxiOO0ytbm72BjVYHGNOD5s1GD6KRQiILieVAQ1Ka0MENer5LSJuLBKotTImJrrq9MxZv
sDov9SmPVMhzMMbxBIdSIW6Z3y0aGRoO2NH8ZuiI3Ae2fBKK0aQb+nANGFUE5k5j0I6CyyjhjN3/
mv2RwpkB0D1VKVd9nqyiSO071d3MLBOHl0FlUu1qFDPmSjldtVBRzaG43lNR6L6gKec7mdCSlfCF
RA2xYedCErrlWjPUXz+T97yPCOG00hqCBv78GPHVePU1p3ccwTXBdvn4Kg37Qu51gox/lPGdncLn
3j/77Tlvx8hg0aHoavpvntswo2WEshLFLO1Kv3mXA89ovRjAyOkRoympuEFwBpy/7M1r8P/5c6KD
AAzQrsPngaA7Yxqz/jKT7MHvMSA+nDki2R/7KeYJSUvjYWqMPlT23HgNrtQa+tjx8N8Zkr8F+uYj
iHrdvYsqxE4bimESKcIMEwDF/yYHmKoPv0mAQ1IENsEFufSCjy8hyYSMXmTmkskn4sb5dZgL6ao5
5HDlL5Z3UA8hbiI/oyY5jHVhoJRfKfPT04Jdd6hapnBnqlgFXsTDTG7bHpuGRqApiJKKGQpx0kLf
fkh0ktgk5hXQEFZG1lTzkP2p4v62+VamCx6AUhUFRzeW5hjxgqf6VDcCZ9nEEosBJ9NamTldQGM4
H9g5md87Z9EKIp3VpBT3PDoDFaTPmK3XDwwfgdQCVG8i35++vFPRf1a4scaCq87KhzWBq3BA/UsS
LP74ZvuCXBgPK0Y8jlNdI7Q+7MAxprhOUfJLhP2DsNqOlEUy7OGHTxmTDwcFbf8hmmIlhPutaKrE
uAm6e/ow0ZTPPSTjtY7sfSD+oLEnjzHb10bKspV/zk0hc2WH68VT/0q+k5VpnSmoDMVJxPq7P5fM
JbHE0+WLD9YiZgFsGGtdaX1Pq/SfIrbMWpFByANy0fqWEuDf4BDoPZ8g8IglzkWmdlwb2mbQ7JVQ
q86YsEjJU3f7R51vwL7JAq0HYkc5/8FIEeI0/s9MujHqIVdP3BjvqBOCiC8ErCuc9gSQK4TyL5yK
KRq5Wg7y6nsQvGZOgJc5JJEy8IGlHIMhQNriPqzYQRHKFhEYrUsk8amSaHIZPlEFc5W7FaOx7Qbe
YxsKj1cAdQ264SYlLyHs77VjJB/9AmaiCYBR+oeFCk93+8KdkH0WSk4SqByIX/EXMWgDGbufK/1e
tFOSJhmJfCZxhbPE+7AS6e2EXjAGPlYBoD9Vw+v8fP7mi3qZ98EGEZe+WdF2oBlasm4OFYNTXUN8
TV27bGkLVuocNIAzUiXu+4NqC7ItDclNByBJYMcgJW2Q5NHl8mpWJPyt8+YfCoDT8FW7v7OILH0p
a+AcALue9756O4I33nppcDVwQ9P3qFkm3jG3OoJglpkluu1+vIjQScWDzxoMzW7HDTxXvAOSMJI5
gkRWhpc3tVTwUSFNSvYfnS/TDVUwggqDHTAKxfgMz4U70pHVA6fbLRNKdl5CJvOSsbcWiw3nqYxc
AmbtXGV3Qi37k0odOntNeZGBqYi77HrsBJ67LER3ufgfc1dyCI4/ZKoVEKpDF8piCZtP4jsxm9Bd
MoA/8BY4Q+NJ4HxW5Yh6a6W9nk5wS1I0C92Ij8deNVT/9l/5rdPtSx14yoZsbjP+aprYHpvF7/F8
24Rx/ZtZEX8xZACYxvmuCHyZ/DqTMyU59VC9oB+Ui45x9T0rTl4BV0xXgylx9JydSxnIkVWLO1hm
f1Vm9rsyxEa+RA9kos+ZVd2lP35uXxcB2VWOc4NbxC06YPGpF+79ZalKqh4Z2kAluURBiigP6pA4
QDqAeM9uPvxFH0Apz2kWvDh/PZ88br3vipHZF3vX2Mpw0kYTa86ZRXDml9B8EI71n2C32jVax4tP
BLDIL3f4pKKoirMnrNkXY7I4ibsl0xqWtujTOdfVLtE1M8Skx82w4o+UwQ8X9m4ImXprUzW4C3XF
sS37d7+bmeOv/gIbx5ZevOBJVeYmvb4THyP+hvE08XMJAmvIRLxY1eg4cJf/zhU5JATZywYkpPyg
t/9Pa8+a+Y1c1d7ufNoiXxz3lUIeaQRAQeTF6Oa9Rw6Nl7T/fbRJjldRjShx0ycJZSTpnn5ZtTsM
ZCdB21vl1tTboE4D63ijoTqp1nRPlnqJsiHdOGEsxOS+H1jTDDfg1Ovqlk9uUXyAHZfdKgudmV11
NZoEHofYAsKi/GGTn4nYLBLjAwHLapT92DdAsY04TSH50xLFuHh3KyZ98BE62LtDARTwNhQaT35I
CislmRZbBgyY7ZS4jWmM6/mt+YyUjsJMe9W+2XnDHZ8SqH3tDWzBy/augW+GPSCV0ET2fp7NvZ29
jUMyg2gzZHInmblgwNTPKuRWF33uxxmRM+g97FPM9/9vPOIUm2rFq8HeeM1PqDGRsopMdKgpyxhG
EWozdsV/vWPZh+2I9d5F1QCp5A9kAOeyBNqep8M/YRQvMWN9D+ourSdsjorfSLAUqPNN4VxAFezJ
X8ojh16zKBe+1jBz5VWI0Fi03D7gpxkxAYfnnLARyNzqpExjJbshI3nbjlO1tT8F4ebMnzYDg1jM
dUstfhm3IADls215jbb88kXGkkt41zzZ7fFzWob6vhXlX4JGTH3DaxFgc8p33/CtbOxIcgRCP6/b
cOi3a4O9nnmnUsyHgAxLwFLOw8lcwb4WPQXsmNRwKvM0yp3eLBSItrlIB+ENpwLro/urkSmMF4Es
KjHvXEF9t66OsQN8N3lF/VAqv88TJUE7c9lbxHPnPoqy+mjcegXVJOp3/KcbPRHOzm8yhMcYLHut
SVeVLj0SZtx0r3m+WKBcV5+alkbIp+nWgeefFSj3B7P/JFnbevq/HbQ7O7AjIst+V8hKp/5iow/T
A0uXLm30JkSKzo4OJ0T5SxjwjE4dYTDD+36oVuLPPrLIE+J8Rl+U+KVXuyFxx1rKmp0DuV5psCxu
iRxzlJwRljyco28Z1nrVbeM6u5r0TagHvM8MmiwKAmcyDZ/beyFUpb0+0AFmt6tv59BwSHZmGlj7
4GJj29XZ223NbLTUwpaJq72INs1W11+IePqS8fZf682VGBOvbrYsiInDnTNmQ0HwG1fRenQXRAA1
L4iuy6dU7JtWYmrnCwPU76lc5xd6IAIvXGn3IjShXMzKwThKdpPpMQZ53ZAM6CRuLrFPUIKbZ2O2
kxCI4Ut0Bdcp53AbLWuYbP+xeQoYnV9ux5qycg4zOyc922EbdCFG0auadcesp4Hj3vHwgBOw5j3U
tHaYAe6qY3sRzx4Oys1FI0AVbpV6TG0D1UfI0Y1l+I8qZoNEsM/KMlpWLVDyBkVQzoKMY11soEbq
qoHSgt3crhdNxoUVa/DWVAs0SK08VocX6haNYzFaCxWFBEbGQs9v7tdg0AxRcPzKp8ZNNOu7dBi2
51fpyVhC9F7ZTLfr4IgBEYvxYMonazeiDAY1khyr7rc4p+nY76qJRhHJbTCfT3M+5nsbbffniapV
QnULYv1Q/5BMx1JT53K0b6Nv2xVdVI8W4u9UHWF1+o42xVNwGZWFF9AsyVVY5RK+jwFTqM30y++H
EpRjcJysYN9TTXZyVjwgUTaQLdJbeqsh7KnYwhQ0HXFzfEi9a9bYvCgcgrkjr5+MvxKAe/2+xLLv
95ZQyEyWqWDFMk41LeENVm7hk7BBmxYvFFZg+uc6lICj+YWas//lUfLuy198PMauR+yysgkKDmqm
kVkQC6xSo6KvJRV6/JNJMw66XXf/zLq+avuhPci71Wk3MRPnZYA/fiJSsiKl/hFjHBHLFmfFE7OY
TbQyqJPg8PAehYzkGRrO4LfLyTeRw6l8vQ5hcoMXLJQmUfLkqxuHvOF8W2IJOMYmJsz6zLoHQbjM
1zZaLBcNdU7F1EEm3eeCynf752T6UNRq/5mC6kwi1rJMLrN8sZdnquHmKnuhdyg4HMxmZ1wSiGLH
mhTU/QKEoo8l9y6hVNhVtKdjRqPcHmkC524suWVc/mwXC3gvXE5e5dmMXe3olfkTcB+QzWqiVyX5
lmazkWHEhBL13+bUg2xllFUmPRuBS3MUouOoOHeuTSwsYNKvdYDIE1ugLEkyPbmmOJ5kOjFvPC6R
EP2Cl2nQnZBq7o8Lb3aQLwjcwICK+t3HY71GCjzNA5S8N2uVKZmN08U/5bGzfWel2/PZmqYFJAXN
0M2Ze1fsxSW33ToKubA4MsRUcNprmPmTA7j5dGWoZLGpN+D3IDDGFLc0QQgYPmQtbbinQ2VAKYxh
ngGfNA7HwY0iNmsOVS1XRrINzPBbTBU0kpJfzBGHhoKhQ73RA505ggyAshBV0VnHf/FjVX0r7ixh
Z5y27j0naMpo5zBIBpPN5N4m1XCNW07l3qdYdr//WgdBBK2h+joh94TA6PYJdVw8lIAEvmyPld2p
GdIhcLWb5QZF5KXko+AVKauTsmlFusjlWHvlEGjU1JYdOykRg2D6GugtmkwqZYlzf3gIcm6mBYpl
CfkkqCtJBxT7WF69fTk9huplTFdM+Oh9RPrqVImxYppmpXQ0bV89KvDT1LzwCqlqq4icr3wQBuwR
7HZVakhdo+EO1GSWKu9ODuEx9aIazrZkoOS5Zd1AoyeUr26kPu2BYNS0n5InZAh3kZgmAdiZjgWa
UV+TzggPXot93VBwfR0MUurGdMnqznoXre5bZNqycUd5pITdlL6bhPUOEPyXQ/gfk13ZhcAMGSzd
cJuxmf/dIZePWybvXF3ft1oHOwMZyZCB4pxbcRpPK0pvsC77e1SpPVgApx8gdKDjgSfQKdTW+9Ms
5Kp0abjV/rOwz1OGQctFnHNyknOYSCKofSFfpkNZdWJzsL/HddjXH87zaOFsLcBiyuiKbQQO1JL+
yCPCMHeIJrqbN6mn21FCf0hLAF31/tEKNFhx6UU/o7y2MDjxh2/IAEhTy6LZY7hCTqaygku+eUWA
rCEG1VqEWwJxkh5WhPAsc7Xip3lwVXJPUFBk9C7YssFjP3DFj7r0ZIufMtWvZ9xhXCsP+Xm79PTS
jW+TDMVyVdkGXWsvGSxt2ZFDDosz5UlCYmfwncR1NC1gEEB2mM5hzR6e2pXutRKR5MUQOonw/GI5
z7Ex17TG/vzvGaEtZjP+r1X0mT0txy0bl5VDAwPK6BPd1zlTpkZAk6ng9wL5pGhzyqgXMze8u3C4
mKFKi/qvceLjxG5JLrRBlRZerDnu0+BAQxMnpoDFBTTc1NR4rN/4p5rwvi0BFtCISjdsohYgKsho
pIFNi83IxCL8JdrDqFZfAsNiCQILcBsbdcyE4wG4xI8FXzZiPIoWchc0I5aILSl2QVr3L9EiXn1q
xzGHAbXzCqjTTtXZZC9P1lH6Eq5iC3ERfLczFq4PwdVf5pJiwxHFObcBCAOJM3V/G/C7WWnJ6srt
F5+LwU3/HhClaRCAew7oevveTBFVf8OD8AodZH9uGYiUYuVhEyjf+1KIBCRkciyosl2W7rAefAJD
gLPbmrp2gyYFwqrXg9OpXq2at0Js1o4BC2dnlVYFdKUd6v+qrNAITrc8L6mhiNy6Zb+7vUcOArXd
xpfz+IRomQ5BEA8WKv5Evi1pL7jrx484HbaGjxaz/bRk/6NaWw1Um4b5v9WjRgKvsOuhLWQ4H2KT
u2YIW9S+vI+h0Kgaj4KzK8dDhVCj2x7HlXd1exFbNlM1zowol4+JGQq1nMYcThB9NmyLEHgUNfWr
JAi/HOQB7VS+QgyV5PX8aC5j+vnzZ4FPlAoeTavhZgFDghyCCvp22BO2vwQrCZMx/M0O209U3Nnk
xfHQUewruWBjzZ2QzppPV7n4ls0Iy6dpKrxO0v8V2R/29+xgH28JBS7EMaPdwiCLlr5txFzquQoB
M/oHqAb1JoE0y9kBbw878MAZH2V4LILSscwBykYYjHvuT2hL5IJLSYGdIe5r2mFkzGGjGN0P9B1B
Zldmngc5BJbXX2hDDni7e6CKyK6E6+sP9XdQaemgWNGaVO1sKYPI0PWOam39DeoAk4g0rhBv97Gs
OPseTkBmrf+KpbVSUCcyrz2AKusi9y71qvuylaOBVoo6DMoTQYV9u0NX8RRematBCDLqD5WJbHuj
qZM8dhonXhc2cVaruoHqS5DvpbUY6jYySqC6NBoy+vnj0Qn54EGuGC/vnxIbvcHgw4TucxuYcxMd
gmZcKViIhRafAYfevtu6X4UJKzRol1ytPZ6JN2MbUQYXhSxZdckPfd6jUVz5MGq7CdLqCgT1K5eI
umLTgyJzHCxRL6XdPsIGLfIIkT9A5AXCzKtfwD2LCqxS4R8QoA5dk+XP+WpRr6DBeaYtSUifn7YA
sGLTEmifBsnGLUIg5ElFYd9usOdtFaRmqmuWwL0bAZah46qRZ7e0oieCf6drP82n5Vr3GehjsXze
Y0espvkFDD8wocFvMnOE5rtgyMif/VaqbI9FUPC9XLUNUCKJbkz/QIuCY5JxpP2rW3ch97VzT7eh
T0QiZNoNBOq9+48a8VNqtdtSpMEX03KYnkelaLgi0yFePDTYrgwH2ldqFP1G20QmZJpE+Ps4Csr2
45S3T2Lt59Wtoipx2ynvnKh1IbRbvHKT9D/G0wAWkzmib7/ZWa7jAhmX73wugKQWFxVoXE6xVvTF
OszJ7H+PxXRvvAcytYqDaX0ZVEWzvQAOBeVD3YjJ/VvoYAWQKIzrdFNtiDt7Y7FCwy4WQDHRvXxU
MeO4AKfrfUTtxQevtxu0SskYPPI7MkyoSwZ4rexr108kGwIvGAG7EgfCKK1jWJLeR9mp/M0LiDtK
KIdBqC1WK5poSg9nN9HcofJq8kDAexYhivf/x1o/zVWlh+deASYoq7onYcG5UAqVu62ZoITXMhbd
sO8QDQdVu6MrXg2QXdoATcN9rZS5S3Ut9UA5KiakWopICT+tMk12kU6AgNPqwc47ZO1KhADWTJw2
M/TavdKJWnsy0rbhh34AwhdQed9eJ7eiJ6s0+ahTJDAlta7XYa3bX5tA3wm9MiMitdE0BF6IRMgk
MWuQykhkidNBn8b3oksxDUUKHIss/eRrX9KfPuanCn+rTe8WLeUrIdw/z0njckFvmGhN/K8G0r5i
OJElshvjhciPnoXGetcDSOx98kpBod7o6PdyzAtSNnxyG3XU/CRaS/wZxs2x//w4A4Yfqt+mxIy/
Yhcsy5MsRKoA2/O4GerE+nBS1NCHXB6n+Vg/c5auq29AmIU47EyAI2FR9hfP04HW1BfIwVBRbPtO
IZAi1hNdGyMdIObg1UvWDUh74BRyqZOClxFhVs2crCpOahsPjIWgvBR+MJ/VNtZP40Pep6yBYaWg
I0RwyIAYVXHAxDgcGFLaQthTIGEQ2wyBRnmpbxLdcBflYO+8iL/MO1J6ggnVHU6/nV9kNyUnR5Q7
fd6BtqKwLvoc1AHpJ5uo55Q6KNbJwFqHKhFR6toYjsStKqotJSzo8a1FqspsOhS8FKyNnNFMJskp
NNNffPon7c6qs1ZAm3Q/VB3LVhG06qNpnjw+As2vXPnOW1tHE1bBqvMI6PhBG22YMefDJBikUJ3x
oUA8R/w5syNzZPX/OMIe2pR4dCs2HZiMdpf5GJ9gkI+hEQCGYfnpgN5zGq5oVKDUGxBWZWW/UvIq
9i+Qvd4QuKLH3HP8uR23ROlieOPIsiPYXfmGWGanRmk4za9J8cYIaF2SQ01WYTxu03wtwBTDmIbv
rVVx48GmZlavD06QvX7/707UdNcfTgG6TXkK5JfEPrZmwBo8rK4nq6DO5cvvX6qV0ASawENEUmDi
ZLInA37uuHz6RNkuRfarCjqtsoU4YrXp04M5eQC9uNiK8fpbwh04jBc77sQ4Qdqy2VNelZ1qsexH
feBwqCvtWB4EMqSxlvDpqUVUaAgtNcdRy7VT0IDk2/CiDG7I/fmmX1OkxE8Kyler2cjczz+MvbDP
Gw6qByVG+PEi4szWWSaRQhKjmAvEkcTtFufK8dBGYW+0jSTAAfOGt3T5RCTkCyko5TVHpAxsM5Nm
tEDIHt0U6JZwtYIQrBluLplQmA2RQD3qEY0I3oMQ2yhbOtQHmA09eZ1N8rfx8rN98+PZywJ1pqVP
Wsh7DHk94aUOsMkUsai5e2YophKN89a/TqHx/duDw888z8RJnQHaOndOhsk00dt2KLUzqFWC85M7
qZ1O6PpQbN1JWim43mMNKpS0DUaKw/q0UMAJcwqLtV356yOWNOxhxC47jsnYPfmOGWFEyapEipOp
HXcbTZk2T6/AkgCILAmCk2n/ycQH+zGWgrkkri0OFk7u4reK6jPSzg2ntk5pnZPBgFoWmwa5xcXT
FzxjuuubaDsgi1dwwjp+kF4PLp9CvB41+QWddAJesmFBg3tR70DGfIp7SFX6eD96gjA+8zaQrI6V
V8psE0aJok0Vpw8B3eGeEiuXSwyyrSHldfhW7t+MIyJowpuh2HSy9SjQzDaWfeC1R84VWlEovfLp
ppQ/UaeybQTaYdMGU/+CusEOO8LLGZdUtx67y5bWd7gOSLmt+Nk9YYx2YlIGe1gg/BEWCl1Y9KZu
knUp6vB7xGyuIrhMgcgiger507ddDeVX8qr1m6P7pDON1GERutrRmjDAB+g6lGY/NyelG4hHBnqz
1HJ9hfkZ5V5uhAp/t8LqdQ5hJfFGsZ+Y1AofnIBXzWnikjK88qsYZTOAp0QAPnvQmi6jhs0dXaTC
jfPLaosN6neZtQu/g+MHOrlz1ekkdwij1xnPNzdIGhc+12IoJfurnefA4aDdrHOTwUX0OeESbwcB
/FBfpTj/yDkCz80YINfgQozfaZ3CTiqgurTWHObPWmuwPN314hXijQ19F5+HoMEwe4kX2D2BRLgx
+qJgFVK5HqTnpQwQZ+xd4FXwlPYuvDWB7iXr5zfZUoMB92MDuiJojKscVjP+WjlRq6ioJyijG11L
hnX8C60VRg6Mefg46QzKnzXVo30aWm7NdFD7cNgdy7Woy71VaFYsmCeNp8jP/IKgLWUvuuhwWMnC
czQtlJdxWC2UqdnfBkm/z/7/6YCSdT2IEsGyHQeU1Jm0xGhep6dJ8SUkRNlXU8i2jTHYGNuVp+MR
tFD7am7ndCyHq0Y0ka1v2VoGJhPBbZrP2W0HzzL8Vu7Qoc7/+Ugh1jPpxm1aLGSTUvFa6gCg3A8Q
BUPRCM8MHsh3TD9UW3M7rpgd1TLkEaS0ARG1jJCc+9Q9psrNNGesOuZ3utlK6CDi3WYwdpZF3kOS
U7cI02xTgdNiiEkTmttXD64SD+bzXitIystcV0PIusGOPZqPZmr0TBZqCKdq1w/fcEmDIQqFA8wd
PHoVitEnBos15zAgcRHUhNU4sKr2bwnFpK1AOslNRsS6JN/9o7tFaiEIqQDPz1WnUqlKMJqTvVda
6zihyuTKBkqbESXXfD/6890UxF9xOnMi41NGvcus+pcNhjl5iNGL8USp6ATvqHybd7S3tO8TB4cF
f/wB8BqoElfzB0QyCQLd0RG5jY+egOpHe+gym/Yf+gxznj+8os/srYM8qlP3bkK6iaQZC7lAcdkJ
s3w8dPBAvyFVITY448TIYp8w+i+M+uSPszt6DeIuRnBCTyQymuDx5SGpv2My6KNwn8whrlxWFeyb
MzG+6ZsYuM+g7xutCy9HrBUNj5AGLxxF7cbJTqk9T1Dd3U/g1cVzjCewcFRwWEu0qwedd4fxlanQ
1l9f0bTROHbak4CXV1yPr6Q1lKtCaT8nz56RO98VrEtB1WaCFijnTYVM6XB0aruR9ZzXxW92wYh6
0CmEoxoI66VJUQPqA6yIoE+wFL1PU83QMg93YAWuwkDDxrEBd77qS7mf0SN++WcYb7E8PFMA203J
EyZ02N5IeVGy1YgNUHCqZvIpFeVxC65Al29BFqAErhrQLf0ryZGzBjlqorkQ7mvJpoClHy7UEBZg
d/+hmMEQBdr5qC2jtVTqNZTiSZMbB9v+sjxZrxB/41YvcrOPEUlJTP1WVkD/ccYzcvSV5f61qGlP
5qAuQOv2FhVW07coaaoGAkqOHLtvGB8VVA7k4KMcO6BWEaHjpxwphQcB6shCoTGQh7ti1BU+ir2f
7CBAJMdmm/SwIW3XKtl/30d5lPvNbknqoeXpzyyPGRxC6E9VHmSNGYGMBR+GvVJ0xWC4SHphUYJ5
0vjrzpZPb2d8JgJZPLY9MvssJ+WZorKgy157VSm8+dYnrfsLcCHlF9z64tvN2d0iK8bYJ6IzrSL/
gU/I+QHIrSXp8ZdxbzT0cn2VAJ0E0gs+w1noR3maXKzuFZ/468euXjyOGHiY1Z9raW/Q4v+ApQ36
TDGRDmGxVk+cd31fuPFxAqOunOofBglfYyEAD+EGm2bTw9dRZvnLg8uZ993HgY7z3SIma8ShN7yw
iHI6APh5jt+MUo2X1r+ZEj39KeTkmB1iDHr1FGJBunwVjmUz0h07La+FkAOJOTpdg8aavGedTq+7
dNOQ7dacKO5Q1h0PmzxlSIaYYZP5fC4z49QRdcIfFY7IDWLQPG+V+BcX9VHCDlcya1ZmT6T6rrKq
LSN43QQJYjLXw/VSVUJQ7Q6eXtjyQtiv40p7Ok+3T/sm5eJwKVBXiR+8wYUQteR6Jww2Nbpbn05f
2F4NKNa6bAmJn2PH7bHIXkp+1KtUsVlEz5uqacR747J8Qn7uUZ1EflUHPIYwdsTUWA54P0Gqpt4s
mVPR2xKDvxigm5ujEnYlM8w1vWvUJz92tFkmfgt1QOk/2ywOx8qRLFNueUuYaj4sGqkgltq05MZ6
k4dEBhNi/VWQ++6bXmBHwcA0ldtf35qiAUJUvWYQ3utk3iXNWOtmgrwRxmiesqZGvKJNfwN8svR+
5F53NXjIzMnmPvL3Im09Y6jimybCykNTbkF/qE5F+03OQB3JVAs6upqDgI4GP8RwSvdw03pFV7BV
1zJJA0WNVFmHSG8+E6HLf7AkVXcNjyWgDoMYT4zmt9TJTaMLkzGMtTg8LT3fwfyn+fKWz4tRLE8i
Yu6yMMaKIHDl9yCIQ9MhUFAdR9vuwCnk1/Gs8Qri8NH82aQevDOkm2eij8KyBhgFmAe7k02PJwV3
sDQ5wULHQA73xVvwhHFkEciO4rQb2YYpuVLMotFpa3cDkQixTavrfh9u+BtrQoj9TzHvK5nkJUQ/
6QLliCF4O4IN0LC8sci3v1XLBp5mipNvepGQBbl+/t9GVwEyMxGthwsmHMRs/seSTse2hQTT3But
77YWesLVXVH/MB4Ccl56H9mZ+k7EP3JPyh2Vj8ttlnrDS8aV5QVGV40mNRCyJaQIe//IwN+XaArQ
vlR6O6AxxLcwK2WCCx6CHyBvu+F9OYNnxrg/rHipLfQ3TEwxarwdGtbbNoLUQ6nUWn+PdfwlGHub
MDr9qTfdXD4sQLYIxr+qucLvgBCnT8WCqNvBFgyHT8sp68s0Zk2HAqocpATwosVkkKJUlkGqwxO4
7sQKvlA4ZE+J1msBFuG0C3gETr4s8IxQ6rCMVzmDZEc+0qLEW4+zR6aYLBM846cvyv8bVgqccLGO
ZW3uIp2K0oFgwFJ5T+mb1E0wEgmFmBt7nUcxqYliZjbj+wVRW9MTP5rvGZ9ZE2UT7o8R2bMZod/p
h8FqvSgw4xulpIV6Qcurc8DfprwTJA42uqaQKq5Hh6CHpHK6aWFi546xSuPoLc92YDtWcaL3FYqC
jXzHdWYjIPpEzyPNBgk7dAVOafGsiFQCXxWDFhGPEnFulzOADIOd5N7i+7ge3ajwyFh3JHyuWcia
BBLou70YI40O1xFxl9FvwekN56izyiQDG4FPDcgwhhFtlnlht2wnMtCNWUZ27W3WB5iguKw8YcpQ
ID0/5HyCkeHVmuqE5JeQ6NgDK+EsNFHZbGPb5BUsMgWxV3f2iCX3JkKR9NNp0fYUW2cDAYbFFAWi
A67NFJ08yftHIbEa8oIJyuQX5nB3qHSnclQ8/zveV/Ys0bGAync8ss7aF/3mHv5WcGP8ETsbnvYk
drEsGIUZcmdHimy7JdYO/eIjEY/JZ6Dn88W9p3O7zGmjIR7mmOQrlPWavQifpSZlBUCJ4WuBar/k
xEaE3KzKnQa7WmbAx470TYrCrfjkuU8ndssi7eZ7KlHdZrckoLMoCFrew6OkUCwawdy9FwFZUmJo
fR661hYBEnfyAPKVFihz7paWWistcERpbt6pDGZo1/Jy/L5LZ4jTuqucKmUkhJntUbW0CcNiy4gS
k09BkkU0pp9esQIms9qTpIdldmhV3P119nDPyMy6hfQwXVHd9a0hJa79I9UfMUQkHy8+kkvq50Fq
jKQgog8KoJI1Ekk6AyC9Vfafc7uCYbOP2lXrRU89fYAB1xg/tpzL23p6aFcV9ZhL4yc1KXiRdbRd
pUKBtZHiX26DvtlkKky0iCQkVr2JMrtjye1m1Vv26b5lFCBu3Nn1uO2OVW/LSIqZtru72MP5AADy
0aU/+AnmcH79816iOBNFiHTq+qdxo56CRyw4tzq0wnQ8spQasdxk/Vl1EFnUAI/TMi29gX1ZSMFR
6XDJO47ZP3cSbewgCQY+C8SOc/OdfFmVWp1z9eh3JwRLhPnYZ2zKyotyJWNjXU2VdAoKUq80KC7o
CL2EMM+8EeEJpi77/T0CEQ2RVQjmZ6CsB5PVCh7o6G87uY6BugA40Jt/JRuom7ZDc3nNrniWnZtX
R1yVJ7l/nMpthFn7tA2OFj3swBvE/Ic34RoYhRfMboZByOiIq6FEjFpTO/GdvdW2O6WnW0VlwkHk
22alE7r/ghxOLGw1P8TygyZ7zBs79mEld4Ny9GQrnrhtX/mFJ/qnWdEaGv1ad5urP+3xkMG73ri6
Bh83jnmKu7MVjOib123wNNc2/8nAyKQMBmpYl9zF891El+KHlMzmNE25T0tovMm4D+6+yR3IgDJQ
qCBa5yYOjGSwfwTZ1CMTFnKQM+RGs3P8bCyYihPk7TTu1JfdseXhgja7Z4hNl8O6C9hYaz89LVpf
W22ZuCKM/CwvPfM31Zoq9Qtp/dSHQSHgWGIfmryGQqq/U5XqT/b9YEa4x9htGkPvqlvqbZgAHb/V
E5HvLBqu74D4DxkLznq/twD9pm5cjW4MZYm66AuLscWz81mXHTCY0rUBaMJYjg1NAF5v3xqJRuDQ
7/E8eL0omqUVmBMdvNNjkiMtLi3BQRnBgsg8oaqLNn7xKXsb1300EitqfiyUcN1aLOo7ANlWvWU6
GeKXhsREmCn3rroDJt046kvHDBdyg1U7DQ32135X0eQY6Ne3V/uDkIetkDOrFmlDMHl5qIsVZ2IC
187nDUy9L8FWJxIRkas0SkXSB8UK+zQJBLpKoG9ns3xbYBjRbx469R2T4wK00O0W2dPUPQoHzkCm
1646KSbCSM5upnYQE/OMkMmXFYk7HqLXaMPQq4ioVQ/kupj65I3a4uAFo6bSuHyKDN4muYO/hU4u
IiSpQNpSKIG5RZIvLtj7bADUNLDe+LiozjBrn/1PULatl1ba8Wp2EFYvISDt5a2rakQg+T4TbD1Y
F1+Zp2gLAiB/h6q/fOWzUZ2aWvjSuW/+wZeMNGSmMZcIsR3rOkP2y9AZGtb6X1VnNKB4AHpg6aXH
TaZDwKh5K9t3nCJKVBNum9seYM8L2Gm1OdN9Sf+ddZwVfp5mRW6gwbsvLJOMu6J9pBhW3gX6ts2T
LT6W3yWQs72iiBYo5hdzeKRtdOn27mSsVT/uVGWBG8T2EtHBzeAZycH3tVpHWVsR9/SVOEIqOYHb
Gjt+LVhWEkuhZienZ98tmarqfhiJiMD0b1q9mYod/3b6Ch6X+HoHpsSEn8gq7oUdqlJXo6RnfmYT
mFPF3MtQzH+76oQkA80vxpLdI3LhbLhw9Ld5q+LUWPoiwjGXHQxDV9dOW+oXgw/DDHoO29rNwb0t
A5qytPEW93h+qnmhk4PQ4le8DnEl4MdRosljhIDH3q0wfX6cEe4JAeh+mrjYj66aS4ypdyolA0IN
0RAVXbtp/5g1u/FuFELPQLKrt8pnZwyC4YIxOcZyw9PhcyaJIxwfNV+aKEH0ScJ8Fdp5QFjF73MM
aJs7K7euTfoDQ4OYQUCJtuGtaJeiJPRGxz24E3EuRwyP7K4RObVhPkUQWwB3nQ4byzQMHyfR9lg/
2PAJiuxdGk1aAD64K5HOtOzo175am2OOmfEPFNMlAIjaYiVpKfd9dJCxIQPjmX3n/yJD75Y2GaPc
y4J06u/KStmzHLMPcuXl1WP9Xs/hOI0DAjZEWPabdC2W+xilDZSzBH3SCSh7pgDJdqPvK4feidMk
gbOCH96yu5yWXleXNOjcfSXZlpMIUMR+3An+JW7I5BeF3a3N0Ww5GyXaRZRGhsk1TeBZrzROxBlD
5veX22w4MTfg5ckzxXYvz/RTLyiWqrJrBn2zL4IhqdPqtRRH104GYqDaY4tljw3do4eZT6hDFT8i
n8J/L59nMupbQcsNE8cbQuguEyKYIuwwDrL9uNMyBE4EfYVQsFD/WuqKAaDFWDWHg78wQrahafVu
EZR6j8Qaj11v29IaywchSmL4xfMxfFNE2V3AiAuc5fOMTfr+cilQo+xROkTP2pNBcSeOXR3+63tw
S+RXPQ0VBref7I7aZuEX8uXguLk14mj2Xkd6kLhvEoM3VrW80oI9ql3ZNwUkxFe4qu4Tbio0EtLg
cA2VfM223Tl4zMu8XsplBjmShge2/UOOAR84v1/83DqgNgfFSXuCYs1Bysbkr3vP16LRCZHQmwxl
wA/Jwkc+Z9OIbeyaK9LlLP071bPZ9s4XPVkVVU2rYILKSytu3ZEK3Z4FRpnofUr+5RFU7NNIiXLu
LAGQSn4gIS0ikONGNO4wU8BS9SDNoZ8vcCR+k2fm7ScCjZtQiKkxRjFQubQQ9uR19EBxkG9qcqxP
8ywJeVURaRfZgmiZHb9GNQb5M2URIhE8Nn79geSYQHbxLJt020hWi2Sc3FIi8cxQTInAAmxJPBV7
wDZZYbO4aGjIQOA6eKevhY1Q+WGapk0fBWbOptr+HF4ZEAUQYXSXk2MR5a+hdDSw1JTjpy7Rz1sm
Hb7qKUcKfR03USR2VtPa1Ii2FICp8oEXsTRd1c8WzyUbmFxf+3rDJsZEEzZ+IZh4KI6Zu+GgnhXK
Scv7nzmdML4esrHNJSxaeAcIBfQmypuIvKZl3Na85udjtF+jfLfwAyQv4zPc/hR5h+9Of4jFhLiU
4wFHLCuOz8ZQ2m870Qr/FdJZgJtCWUlcnxU/GMVN61wH/TQZDig+PRrjfl8xamm2xHIsr69s3bAW
lGaZrMh0uigi3pasMSmg7Ltl4IFka80v0772kEmUWklMxpJ0x98UtQq9VScEXRABvDPCtq24qB0N
enBeuYUNXWOtBwBYDb8075sHpeNyGQwW4b3OR+27JE08S8GnC+SK+oaxR8Dhr8I1Ef6IUsPEKaW7
XG/fA8jUR903I48UKjC5wy5NutGzPLAdLIh003cwSkfIHG634MsMAYiggqFvLXSO/zE13jNxSS0I
QFwopu10GmQ+6xSac33Z6yS83WO2ej2UI5d+Bmbw+ZWv9Y3ZIWufyLgBgkLTRTwP0xDOpDXo4KZA
YObVB2p1CnKlp4KHNSDL3mu6f1gayDHM9511dZ9BcZ/kKEb6n3hfikjpX3AKstIGsvKAoIhTZ0Uo
Vfl5mq/LvpKCYwBCLGEVKecRQx9e77D35CLlXKQgKct1Yw4k2MsS0kd7LWPkZN9+8EjpaBJP2GL1
kGWZUEVEIbiDOnZ38I3h/ZfMTYVx2EtUTUvHp2gwT3JY3v898psRc+BvffU1R3cEIv2wF/fKrVrH
hvSjgacc4rr1HxkXwJZSVJqpuFRqlfFgdukD4zl0kSFDEZ2HB9aLyiqqgEr4CO+5WNwtUaG50mAb
h8QiQctOBM9qDFzU0drZqU3wWIQGv4WsJ2rjOJcNGxn52UToTCbPQgFVDORpNiOJI78iDQQMDy5+
UwuLyGdkO7IvA8I2gF36WSr0r0WWhvhGPwheheg3R2z7RRnzgaLhTT+EDdRih2OQhQeNux1iBUOw
ILokjQM3TaZB4YpwZ8scNHtAEObcy7iNuF4qSkpXsBFqKDcqDlG20lD+hDWpd1uJ09FmsHQ0/h3l
T/HFMteww/p0YbNjRxDtY/1DGM5NsMwBpXZhLjzlA3dDnBhhiUeoFCJMTC+0iU8t5YCP3sdLqRQ3
Z7VihI29db4kpxyzw5vlfrausbT9QiIc1neE1M2nAVrd+/qILL1yW/HNelkog0bb/RqV07gtklmY
dLLwo88isoGRXyV2c+EH/s2K73Mj/aOBaCbGyD7rqVIofT1LojmdYsaY2LEhvUueMvkzBO+M4t7o
mBJsMt6jlR1QgaLsgnhd3eDAEzLmzZreIDXAslSnExLpXek+8pFPL2HuXk4qq1i0SLdogl/147yf
5qRC+1zwrq7FQiF59ISKzUMDstI+bGMA4jnj9+CcakXsWRxiO/ezBdNpUhZS9os1hNipzxLtlb3G
9BySNf8zMSFpt+RtwMf3zMETJSVi57Z8+l5Nyf+toOsnwHo+b9f4KF4jSTXb+TOL530ckL+ltehO
ii8QuOHJGl9tS5t5zdacoRAYIo1BLcBaCgiS0H2zdGXy9IxyPk5bHxuyN8C9ac4FtgTnvC04fHao
nvzc9+5DfLKaPoPvg9WUPmF0H9PTuP4k5LR6pjNYzay2bhZv93qTsO2+Trr25m0OyOSJ/blwVY+S
tZFKDGS3IdG/5dIZldkXoXvVV0NIF6DLBXh9jvOvNqeGILaflQK+fI81mvo/rqzDQuzVBc9CypoG
176qB6Iw4SRQzM+d3Q9Eo+5OPs/fU3K2vDKeCcF7cZXtchlLW8ayoPfExw2vH53yrXtiKSdpg212
yP6fRlm8sc088rKK0c5xXVOVaCvuYog2EyFRJlMlx1gmEGGbUD4by8WxbH67NYa9e7vzSmEJV+S1
lkGDNDinOY5BSF1pX7EMDLBd9m+aAkG037s8/MgWcz1rQxd75j1JkXodu0QOza2BHRUDwgvnexFA
gkCrufQ1TLTUsrTkbWYGSvhguQRmhmx2NE3s5VQIN9FyTCyYgLM0Y9SPdWkLBGmJ+3nPmjJBMlwS
8z7IU76+Gmj4aNdWnp5UNq9Lmvon0QTbFnEjcgF8SRdBHqGAdVSGGkh3vWX+abXTBnPw1jXQhBAg
nkW5t8CKI6kNtCWKR1xQ6eJBuXhCcdng0kvPgZNLmtZGM4ZATGiCJPrQyNa98m1Ts/ctLQIy98HX
mpnrhzXNNKe09iiP8qH01P29gXNAu5qA3GzQ5F0YJIs3vWE71MFxCvEnObtA/+dZ/NnA7vTeiJlM
Vwf3OEUZTTAtBc/7DKseh3x6cmukaJHk6FKBv2ywCo/KLK1nLUIZh9SG5tN3va/U42bsNTKZshLa
J/a1SwkYYT6O2TRA25nh9k7mJnhfKWZwEZAuUasfvw0Uw39VNDk6v4enN6Mhbxy93iXp3X8iVLDE
NWJEpvTzXD1sFsrZ13MN/R1jNoYYJ09q+wiFbvcB8egq/oAb6lfUvU35qQi/cM4ZRmu/51EAVVpk
lkaZiNfuFi4763K3jnx+Vu/rmJLZufgZu1hnZ66iDpkDCBbhQgCpQS4ooF/2hUzpqFzLBCW7a65m
o0FTCYOEkECsjTGlMyQuf9XW/lAhfnEiY27V0r1LVlz2o3SiAdiYLcfsdCWYwNuE5rJhFHhFCyUe
gpUWshCgnI/9XD+oDG+Vd76tyr2A0kmAyI/93By/mS7TU+rhHTcLl4SUJRMamQDZRZwt0PULkUrk
Xwo5EZG/SVtnnO8dXFWQ/xQucB8MAhKxEajHRSxjgEga5RPFvhQ3vdyZJMBfH82nPr0aFKQJC1bO
u9SG43kFkQ41QiCWaT9iei5zqEHJtOGiqoONXG2/7a/NEEOgmhHB7AsIL0c3KxyPUzkDSRvBEcHZ
CijSpkyoAPFx54qawo0IJmANU516UWxomfJFyZPWvkhEHKMMAv9XyHWPaV/LRvYZ1f6xkbtNN6NA
q2y/zzkziXXOfLzcXZFeM5JzA2L6iXXD4oba97E2JjVxo3VL67Ttk/9RNngFoZHL29nDy54h1ek3
8cc1GzVyeGGMGniABy4/sNsDZxS4E5dS/Z2eIB1f4e5Kf9PgawzILp6yZn3tMMn6PqXmWfv4GYqD
GopdbIEYtyghYO8KjDSaR+/9/mXG3OJ/RGCKTQQnEq8MZ9BCEg+UWJxZqz7kwGZd5wpvFGxUJTNA
MkvsJT8FZF/B9QWv2yrnSyZQWPYRtAjzPxm77/0e0WBGXXBt8YhT2Q6pyVJ2vPTk/QyKenGtFMeb
txJiid1U2EF1l5lggA/lJTR4w1KgyTOFSqqZEEihM9W32bD7ZZ7r6VDAjwLdNASIvTJCzK6WWXR3
VDPNqmexB10qtDLz8X11kTE4v3EQU6M9iZh73x5vewkjomLkF5QE4CFpz4vISE5CQpX3CqMbwRnN
4yG+bbAyXqI6Cvfpjrsr9Qwi1BTHWgG+hdDuYxdJiNrODfVMxbMSeQyrw+nrpT8eGS8mpnMC/Yjt
EjDGRkMcW8ceQi4f2PB1O7th6FF4AC0syfXjJi0VCO5/1mCIkqqnthfC8aT3dHiHq5VNnhsI0j0F
K3HDiw6MaM1SY7lyE30Bn7kf9uWmYDETWzxak5+82PVv8h3cIXk6gDpGqDFmoSAYKYHm0g7auQhf
yLeJWoqZxHM/HwGewoff9c/DpC4iV304fpoiRNNQiypTcz6fzNWHy5Jr6zX1Qb5vJ3C38MHM9Vfz
/d5IC2I+fFkYhb8NijdEkn+o/xc4bHaAkciyD3OOlDcHz5WeQxy4Ak5EFjCQxVny8ix0EAA/Fkuu
I0bKGS+fqpleW/RHXN/eFc6GtEQ9Eq7zKysXJFwtiS8fyCYR2N8tYr1fGUtFw/kdXM9fcrrJwTll
miiU36uXmslabWBMqUdo8xZ2Zy1eM25FwAbxDaAKOmP/R+EHnTLfr2usj5rkF5Qifx/hE9kVhdO1
IWxJffblY/NlRCeZMwtHHyLSEBBdpCmBv1rj/Vt04nojUrOSQ/YwFrEms26s/8vwHdYIW6ZleRdJ
GCdRGmWzRVKjC9cilYdM75x7R8rU+NtCBFmCQd0jU9WJyEHGCWmVsCOldGNr1a+Jxkd4PBKogii+
W6arWgmliEc7XTxyiTSZJNFEXHumx2KvBxedBokzRL6FLBJL3Y+0c6tHVbm6VBAlYh6jKoK7cgm8
+CGDomYwKine+nAHZVP7OgKMx7dh7jxUl1XqjzwqlZQ48pEDPZQBDIvb2rvd0ECQFOmZ9iZxXORM
hZhUILEqfiTqdP0I4/C7d8vv/3rgNCfvYLzm4lonMJE5tpCDsKQhNogVupdOMdxzpSXuueJQOIcI
+S4QUk1GthE3cu4J8ycOAD0EUJolTc5Y4Hi21lgPK+EC3zqLLgOLlc/og7EtowNL8MtJm+LYU9fk
TiUkL46RwIIu+CpfCO7d0Rm3eScXcUEWk6wfP+S0LdfHibU1Gi+39R87pywH05heOaNVwoyQvgr/
MFGY4aMd4IADaeGEho02zLcujEwQ4gTG5MSyDqjcZUdqRFH+znlstmtkL4v7fgEoO89QvNNajfZs
Tsvk0H9o60pYRhuj7J15k8DXOsuFqneTPwPrgH6n41K3svySqgPqKb9ZQRpjPX3wX1WUk1oTj7/M
HyqXi1OJ5GpoPLazjZcyl+8ds/sMfHiiPt+MuxZQ+QybaE8rTgPDAJZHhbhQ7/S9D8jMVM6lS+ik
ZGy3+MqAu7vaH5uCuwqQLrXLua4Q++6GpqgZmYxwPfPNeM7d/MvltIhbQtjS9pSv4gQ6Wigl4i8Z
NMfcCn7929yhqLKCfyU9jyPh/TvG3xhPMg07pFlxxAHsIC8OBfDoEd9oTbl2kBGcA5IV8XOT+m2K
wD4ijryPz/riLfqmyoZ19SpJPilLmeskF/b8aq5DC/MU/u0gX3JmJJpI1FGMpP5tTCtqjkaciIfA
oGQIGkAjdeyZcuw/y8d7S5vtdvdQa7XMm742xSeRU2KGMt2mzQqpvspstngPm+J7yOHhk+VNuCBE
7WzELsYxhnAMLEBMeiIWxQzGOVC09NVh2gzp/KWqT8q3zRTd8OC3EG3FUWNqXMUzjSLBHVaU+Qqj
uRZ82NYy5/LGyB2BYE01l+59ebDS7XPGl/m1G/hF8l8twAMwhbwEjuR4reevNnC1SZ1QE5RNhqy3
GCCKE/tHAHOtzGH12N0gFT2n7Nu3nk58HZTuuN7vMBmx/nphiVnUEnibrFaHsmxJQpajJ1+nzau4
02CTq41kZUVFEdqslPAb4dgGgUvFIyVJSfgT3ig0/wnQbwD6SFSEnUCHUDfxNnDO0iFfLsb9qAC3
INgFl+wkYm2XQPudm7O84OJeHMvwnOJ5D0ibDOXXnVGDw1DvrqE1b/NxLM7PTHmDR3NJPCoUrlf8
677pc4NrCtk8cNoJJWYKxuAMjZJ3X9BSiLWOclqRSC10UI7BEJ72dmTHybEzEZG/kmURdgH3vzwv
fxjB0BhD4DxQ9oorgSheVmdrspbFBkLu8qzjRgmmwx5WbcAoDyuJYzFDGnH0txbhCadd0B7st5vI
Xs3syho2ZsHvGfbTuQb2opIVbuZCmmB5THWQi9jpEUXhpLicvg0aWhr4bk8OKrdpaV1QcTHFJlvz
898hVFVjAnhcxDOQQt4i53N273GI2yl9LDayYNLyY2J1uZ4sC9RNtCGsVWpaDo+Zmw+hi6WvWv0O
a1vslcGVTUwkSpoUIW1V/nv/AwfZQHdmGKeZSWqYPd/Q9F5NnlEPH9/ovlhztBA6i/5zUPNPHJ5j
YWjV/hgO+zifJepb74xhXoy4Bo3oxgeeVvXAvKvZMsacq8opGDN5+lv6eYnhF8OYPBjBSJpp0dI7
e2EjiM1cU2giuAu2Q0zugW3BHc2iYDjWdgcl5Pdpnqe3/YiXai6wu3XGuKTeOJSi3ZdMFi5FoqnM
JschvPd0h4ovq7iXEyE3OZxAaMmAXUiwAqPBi6AH5P4D5ST5kJYyuhtUQ926mA3we+fEna30lUdo
Y8z7Ip9gO6vM7ZkSrkb8PtVbHnyAjcWcwUkC6fOKf05RPWDBdAyaQIqtRGPwUWkjui8VhSbzWhNR
Zr6k0EeiKBioZlOy9Tq4QpipYJsdpnSwBkN3A7htWl7EY8wfWZPmXCCR5zucnl3IC0YTQsq4LhTE
OEqSOSiGxHxrI47Ydx7eSaOWFpkqRuLj4JFF5Dbkp/CZDusn7maiBtZBt1ZJZgpzO9+XGhjn8uLo
HMoYn51RDTl64lQKfb0XvWkCWyKFAcPo8n0XpRAkXjv11WPwqPcJI14eLlobJxpz2ugWL/xSwMZj
Mq/vn2BXcGSZuF/OhiakbbOZqZGjnIiKVITlMZbzIsFfo5AilCQT+1fLLICpOelUXaFB7mH41tlj
I/ofpjJEs73+EQU2ui8TZoCpIdGF74qSnF/v9FTGBkPmhEn15raQCI42SGMs2fA9tmjrRB85fzwH
GMhLW8KgKPPLJIpKkIJswxUwKEfyaLJ4e9sHuJQaJNfI6NJ0pCydHCJGvg6ypTRKf2RbOk8JooLe
O1UyF0Gx/9Dhc/EV4zOltsXjS8L3qnNLOEAh7rCnAuagFTV81FZJR1NOSl/jfJR+k6hXSBL6vJYS
wMZWYMVS3jfkgGLhYzwIz618Xmn4fttZovBZ8fS+ALdjo9FjS/jVG733RfibOz41k7lr0WBNG40q
8+q1zNPAVa4p41zzHgVMy9ttjlbnDb59e55gpvhxV+rejQmW7iBdlxI8j6ObASKsmcreISDWlnew
fQtULWfm+Gaw2zhTy4v9WtrLRjCPhJKeYub5cVgcwagHh4Yxf7ywGzyl64CriWhv9kx81RMAG0KF
S/mdp7B2AXzgUvHJRsW1g4kHzmqSTY9n9nQvtZhw0JSrKqM4TxrZPNCIr0iAxO9++V4F50Bem6mO
QCnlng5lTbbiHYPfQqBt6P7aKx3HkvtgqPvrCbu1fJHQ89XSyWJfCJVW9NAB/pPo2N3ABzW7MFCE
AmD/Q6nSLuQUy9LIppuGs5knHjnG169QySMg8cZ5GoJgliUrIhIE4CIh65M4huvEwj5WZl2acWk0
EUZ8BgOMVasCRhusbD1WfIRnstNy8btqwSBV+ZNQro0cBuAUxJeDuy1lPXcWeP8iioQaGxv6jorQ
bneQp8M2+nHQRAE/X2xAKjwM5uNrqV6f60IzxzsMRLI4+8ROF6GgdMiX93yLABGbeyKVpDQ7TqrJ
kxQfJc2B0faPA8bU/0pwEgRrtmDyFYP0aW6+LGJjQXDNgL0gRmceol1iROCDUURKNgrVepPF2xCr
t147gYgouZyAAB5+9P07FABZZUOt7TpteGCpUG88gpvldu2l58f108k+4a9QY/dTFoVr/5f8SU7O
FAIHLswF+0Z9kGDCe1Rpo/d79qAIpidx5ERWLQRDEDbPlTnZzojCsUe92iX+4O+EppZxjptTdPO0
85Y6cQV5pfMx3N7/xpYCV4buSd8tYRFXSQ5Fne6dCTF5ViHqdghqlot9NwkvpzgwNKiKBpWCczmJ
XaYigg8cD0CeWBeWt15/vi08uCtgVvGc8aMbsUAbpzK/sLHM2q9gbeCUspLOPivG1rpzL4womTiR
HRRRSRzQuIEXS9++4UE86dp2QRc3cQMXfO6mMlM9mBN0i3nXaXcsjJBMt5yqEOSgdTnQT7Z53q53
fMiFanRno5EjNh2Vbr/xCbEUe1rJ/R06kKMaYnwwFKkWaWXNcp0Pz1dtfmDbzE9B5teyPpmf7UhD
pHq0LIWq5cWv6l/+j4Pd3euMmMVBPd4HziECckXZwjsiClBHHmYB0CR7f6bLJ9ucEJV0nQTcbSpD
jR8J4QmpdMn0A6Nkh31D/Hs4cyaRk/BLALwuOq+2W1PW4uh5GyQ4MtQ6f/KM267vHNRjdPwum+9i
dczqm3GlVtduoXvKOoyFmgs9LlrJTk5XIOHLyPl8eOC2i6824G3TMdGNVDKsxVQT98HkeqT8NP9P
gH0prT6HxKYyGfG6HeT9aoDqZY/rP+WlP7fRoONLFdf2UaZCOaK5prvOzC7ipUqLqhqMpgT5vi//
UgyzFnSxn3Wq2EO6fAA6o5cUocKeQSRFxBg4sA0NfnkNmJ9s8QNGHDrLcikQkyH053FjK28/4WcI
TZC8h1Z9SC+8noCJT5Hxc/aVNKH0xLWzK07037tSPTysn+S8FP2GLZ+odcJlBhvAWFDFevc56q7c
52JrEQLkG/DvMqKFtrmJcYVe/vrKPxCmRJu2QpYNHdqc0FCDSCgSyeDlMJhZBzYsRe21m9d5dUJ1
4SgSpT5ohpayPQnZtFNXMP4ES+L0pxI09qvcFO+cNFcIWB2yvpIfZ46AOp+IJyUs6BUKWuxZ17WK
egK8SsguopCJIzvErgt7lTclbmFT8UoJ2YmmHvoqyNQC4XVdqU8rQfZvgX00zz43TWgDqXsmUXv0
ZA6hFoNqTM3wNGyiHTAgZeL06FZIYtSppih+yXjDNRiFvJOxnrRG+lNozdZl/CN2NDYdPSzACKai
7/jjnpyXri8p+CBHwyRMOnqJIdF+EZTZ+ry/Qu3Q66AFQkrtq+1WHtm1hvVs70/gAXgjvW2MHVjL
vFMOtgPJZA8S1vg3L7dohyYPIQHDxH5wIYAiVfZyQmFfT3rr47WHuNRik8iBE5Lwdi9G/GJgW+/W
qSZUNf1wkpIrfeSSlnBnh3OMg+Fq0TrEWW1KGy0Sn6O26wKX9fKTswAE0+BCQ+/ZzgrHMPBd9aBi
5RrMcuSRpaO6QW+K2CKjE/wLQQ+QHfXT+tcKQjn6e1soBIyfyMLFoGJc9VJ46jJJ/jKODafzxWiX
si7To7C3JHH/ApgtOAPbWcuz/ij+KKuegyZ2Ldn3j5pV09eagao1WxwRVcCYx245dWLxaLJR+x5o
PX2LIPtkdSMktQNwMTtsCaglrwkn7Qk9N5VXpDfgbkSVuvOAgLOCAXD9A8Stb5FdTt7DuThpij8c
6SdOjQnF6Xphdv0WeflQjcC3BNCnKRHmjtKxRATFo78X8Tl79u5tSxHARHQSgRn8hzbdYSNJB3as
qBNvDu+wktFShHbDmvcjFRlgHH8rZhmJ52A0DrlA0sh1ZjEaH5pL2nAznUErdArvjSkIvEWknugN
EMejyhQmD77YNP+C2IVyHt/SSVhrcKUCevD5nUQF3xszfEXSlPvCxDsqeuMZULgPOF/ETf78h7Ob
dmoC8wsIjfluumzJSh5afra0jy5mez/GHL7PdOhDIpG2PjXQGTHQ3rhurcUuzw6U/GeobmjNLOz/
dqzprPYLvnJ+VKi7slhglVVzs0IRcyDkLlCrT7XtYIG9VaIVYJE73gp7+BWGvAy4QK6jj2SYKwFS
SjoZV4JzkRIq2OBU+1t6CVQu0nm5neQiKdw73FdjOF0Lm/aH+WeKogeDkzDbtjaSYdsVsEABbQWW
tAz9neryummINnASrGP1lJW3m4S1TIRWqB2iuzHfnQ/RoYzEwqfA+yntkQ31c4cWi8i7EVtDyh76
zbld3+hNp0IICgCv45sXL28B2yKQjnZ+lFuXz/Y9cJ/FdtgvDpweyAiMUycjfeYsKvmoDc5xZ/Cf
dqRNzq1bXBRQlzjicjyQx+w5w/+ss/RoOWP9CZ3hnKw/DgbYgIf1vc5MgoMLVM3cVNLF5m8xtOy5
kDCORuCJXvg29B/QjxDeqGaGSZeKUdHXdFr4YQ27O7Q7JAsXO/WyuBZZtR3/5cwDIDYlCtg5TJME
j4Oe6KRgESYee+6T+Ecxep6IysD7bKIw1XBEj805O8vLva5jUM4dzjLAFcwcsvq1W6VGclO3JaY/
wuaQjEsL+M+jLjKEpR8j+jtbX5AJs4/9+e7iMa3GCIWGd4bB2MvLgcB6iISYzy2t+c+aS1FXoSF1
oJOUJILXLUYq1xdbg+TQic0V34dsHyAvQ3TTR+Hy4oEwNTDOjo2+ARQVMjunNq1oOzlKj1lN0jaV
33BVJloYTn551eRGA0Orz556Vyizu7u6PcSk8Ndam1RkF5OwjMvv6ywoxefBgM2rzXYrHq8dUlv1
bxMgBif6KdZV1Pwe7KIFd1f5/xC68WhiYmngrliuJs6QizabIsUxh079bc3SHEQ9f2Q14dBYG+9N
heA9FlSon5cridMGVfuckuf/itulNZEqcPJ8hsLDwIXnIl3/EpLU/sm45SA5eS0H9mHg/+rPB2a8
AEndOU25ab63hEXr0PqXX1glF8VTfssGHVbXRlBtbFRQe3XJ3xUXBft0DdDh2Ma3gv+RHKwoKhhP
ox7LAnCuDwIXmJI/C+rAZWp4gKUMkd3CEF/y2sy5Prq156CZWRwLIcx8NE1OUX1MKy5DVeOVd3lp
BcZj2Da5kpwFWu5rX+8cAfuyl+nlFsc+xSMbAqNUPRMjEcw8nMiVELIf77meKRyLkFeTuPRlG64F
nTWrG3BS47vQlErb7i0n4LVvCZ/Gvf05fWN2JVr1a9vksfIty4xMVTmL71P6VFNOpcFJRVENEg+a
9sHbvgT1uhvjMRQ4a5JE7A5F0R5+2G8Nxw2r8ehjw7etT1S1UWgzt5S+h6xgflbaeROf7Q5eWwea
NDMbEFYAXJINS9IJVCtoBQvZvahJjaGfPHOu7TqcaMAFK5YU8y4kfVzSB5yk+SKFM5A7kr7Vk7j7
vMktXlo7+P5De2P/uQXAG2g2cnqyM0rZlxvil6ckQmqZGkd3LIq4BxTAbk3f07Cym9DO7SkBUOd+
7qaBSISEoIciwTBuUPoLmoLl5EOJ30+yE4p04FQg8RQyfXeL5KJcZycp7KAVzNpFC8JbL50M8JuQ
mA2jSBwG4P5TvAivbNkPo6R1zAsJ/rJB+j0lIpgyEeJMITileROM0Y23CDmYeTSUJhNB5ppbhbn/
GWb4qAjRPwIk6TXGSdpOonVANiLfykj4V/Ek2RDqIJubGtygWkVdhQq+X2dS3vGd+xrIbNw0ypjf
1YLXYhlZ+BiVo/3pnmVOtz+GreIaYrIc4cRqUedyTXfkR3qfd90DRJllU+5zOEkq7BoXP4fLz3s5
Wera5gOQlqGoHpH+kiImsvQKIIxGliCZvoYRtw60I9yMx02WoWpqvNgyP8Km2ZCqkuxUFSlbg/wO
AX5kl+zIRrHUEPYtrl6JYVIKgQvkEEgA4kKWUSCq6vy2oYhIWcBHmBLMpRYQtDo9gqkmBQz45nOU
ZwazfE4eSUcjIogeqO+2xXJyIm1hIQGxXsffybhQvRXBHchCTWPQcctCzGFrPspZ4J/W16xZIqQH
ZR5EUoPs+/7dHb5rFJuwi16qQIZ/HMfFB4DqftOUWvTtY4uV1cdwYWVY2tQX5LGjzrkhD/QD/AMJ
m9z2VIhlaHfXpd7l7CY0hrR0anbEoLy+wSmD2imTS/MCo5yp79XXqcjL6TGaXNK6vOV9XZslbGc2
3A3FsxRNDKk5ZfKajO2yVxU8ANv79m3X7dz1lKkYC+cvNOWetvuQu+iRXwnvJg1wQSE0OysPw+8Z
C4NSnqCSaCek0BNVBQktrt7mr4jFb7y3E4v+OHhW9d6MdJWbsa0+F2zwv+08VqjzMYCuSZV53DeC
fxWuN/JInGNnFE2C5vXxaU+AsfehwEH5oLYDnxZyUzfjxXVaUyGAk3yG3e19Tqbn5QwOPLg1W4Jy
4nebwooM/i5y/A+OxdNNa8ouN4CtKD3hzWYqFUzZJW9AKqRMW24FWn+RlLDPSIv/0gA12Hab1YE3
toVSxq3y5tvP7k0JLSfqI+/di6XRm48ZdRrUlbBXjVXGyhEqtpU+d1WQv59ySuW/C5Sl8Qw88R4k
opUfZyrHhDZcCKz0BinNW578QIJAdxCz9f/DAe4aCRIlh7k8j30/SpT9UlXit5tM1FrMPYZIalWr
P/PtCV57v/cPx6z0wRIQL/qMi9TJ0xcS6u2GsgS05k6gwuSO43EIWqPaxPcziLgs+LEWgh+1eSMR
RAMe4KsAdt6BWUNxVhBLZ8d12zvDvnZB8/e4KM6KVjaLNTEx8f/61al7fPWCuKZsWGtDMgSaXU9D
7EjKzFdtG+WJjTJ/P8sluJtcBm8Cz4R2vdj38cDgKDxPCJ5r47xUcyH3kCg69E4nPH5A+ZMxog5Q
5BtBATCb8XjP4V6VG7VeRf4XGSmh7zIIfXR3oExeCZjslQBS4TB4hNCDVmto1MMKOly9A7pWLxJR
oXINVSmi0mCTugrfKicGBksvTAaypMFol/kipGxiF67Q0/CH9tclGbUb8HVRvdrVNmJURJ5yWzWM
v1uknF0NVa0nhQ6hT//v31nTHFTnrgFQd0A+45lx5HciIpcN7BJyR5y2kKPY0bSgraU5pfjqVW91
eHd/bQFhXIVxvFPlAKeXseaWZzpf0abaRE6D516oAL2AvnO9smYbUtPEVxhhK5mW60iZBcpzQs7/
D/L9aZ0gQbHZm/xsEUtX89txoSS0yP+cmOfIq0MetE7w/LWCiM/xAdAtOZqgDOmj4zGdmnexIdS8
29Nkw/vCDNP0LaL8a4BciGhZIP0QNhHgPGRlC4WuGki86f/Un45eWIEMZBUD0pLiBBzDAfYP1ZlM
w5ca92SaPBWqb6ShxhE+mExg9I8+ecye5SY767RcbHc/gdSNY6/zpRTb0PE/uDURZls4Y6w0o8mp
xHVqp4qzJwMiQXKnnZLwYA06ZN/EKcvuIfxIPi2n6C9DBJ9bCCBrQEG2OYwqdgsR8+ZqjCV3ht96
dRE1ES6ggv7kCwpd0LoK1Cjfip+WRMZrKGog6+aFkdwpuABj3K18V2ZKq4XOMRyL6tWE+MutDPOT
6kIPEjr+ud5WEEG6X2T7obJueFb4AT1oQ+FWRJO+mdlkP00E0VW4Dh24N+egYHV1STawbApv/vdj
1yQmtAuyvj0qZKGejwLCIf4wN949O5V9X/dRAhQgTkBoYey3/PSA04azkZmQesYo5Fbpfr86PogB
4OJH0y3lVN+yFgO4T04fDF5ElsbEbUJiuV+QE3wzhyh6cBB0f9cQotX90g7lXQZi1PEk1TFRrnyE
PFZ7xtc90dmEee34c6FHZWaDKOWnoMJZvDhTHDO+fIATcfHbgX3S3UvEV7xfRYcTY7hqpfBGMEDX
Lab8jgr8ue5slIi8cpRxpAy6Oo98/kBqgBQTPR9ZRS4KVL7eFmJzQAwT8vtwA21O42qAmRyJY1DH
UCr0hbRebzOgVCcWRMQNVCX5SVt4tTFpcDwRRiWahL6/jVe2YUsAFP3jqGlJ6zG2GD3Xk9u8pO7K
OZjxTnrebOU53mtRua/MFrbCEaH8cnAAZDESxFJ1QTDx5nZGivdQxvei3pwgzGalqzw1Qwr8QVcv
2E3NxHz6yd/jKU/GPR5mNJlEogcuxcqO0VoIFiwgVGRRX6xDtTqBqUxC7RBeocYdI86Dm8gWaRAO
xvkvqJaGyt9ioQ0Rg26FGV1nSfjmAKXy7Vom4a6QEmz4z+15jb6I3j/1caqO/zY/YsXbbwH/h6te
FWDQf4aqRxa4EiS+FbRrwGvu47c7bjzdEASQT6HqTCWkCn9Fr48h54hjoXYqQxx2u4UG11TwX8SP
k29I+XjMHwkbmm3R+1o+khvJYUCNUkA5xgUEosgrtJLAWUr9LElgo3fU+J+qNa7c7R8j5acX7kAX
holzLbaGQKCReX1MnYbFWtecIthsgk7/K8dl0Ux49ytbFO0SgaqkFyAgyZhRYXtpHNf3YoxgqzXN
j5Do9zr4aoifmpBKObJnhYnrMyJ+76KbUqHWo2/5DM8m3pkATWVQ5pxdTIsvbMyyS8o/BMZCSqe1
bhAU+3W39sY1wC6OkQVPjxv4wRhuTSSGS6kaYv4qTpylUZCc3vBYB/mZzUhAo+kuPD2zkpDybsUV
nFVmeEbwY8IgRyHY0anXq6yuzfJJ/eRPyvm6M+99+Hd1F3Naq3Eaquf7xWg+amy+u8SHWawaU54p
7X1+ZjCNTsfwtGHX0VaKi3rjN7dNRX6HpqFztTksHvcNezGbcHiyTT9CcrPVM1BQrA7HLy61jwPa
fBGgbJRCYwx6IXBvmBJeQTaiHW7lPWh7QOVrOXtegL/s3fcWhywfy0OTRS3S1TORcql8Ay7GU0iy
36m8rfT+vXgsT0ZS95KX+eqWgFMp61Qoa05YhoyO03BiMPutOrvgFVAWwzcfDwoCJ60eR8sipLrz
I6EbbT34mSRQpS9Lac5vAufMz9rH0Ktwf8tm7gnV7G0cR/lykvx3iLNQFUeaaXBlO97qaB03Tj4o
+CT9p5XHyynRynJ+OgO+pEBypG/EsruP5hShLT7i0RMrZZnSEaJ0bbmdkSZhw9nlbTBIwdkGe1BE
jGtctRYMo3S89Bv5yeipMnLj8pKPtTn32w5+ZtWVYrX9648wMcQYz8V/W4+vwxTnOYuWJRI6WNbv
cNuHFMu3epC220Ikjny9pt1rZqfAW78Wg5sl/JzFOmRkijNyt2VA8yoUTjvOemjS31EOrMxNzdo1
cQNSLW+oCiBOSXxv56/7H+30pkLrIDLPr2PT22zRmD4E/t2qSN4VfUnV9P2h4Z6XcCSeIjBIOlHV
I6P8XwI9+a6Z9yFFM6mixQNAitPDPu5S+yuaylZ+uKeKNdqSraFjRn+e2kkPwQDFAO3bUdeIeke8
QA9Kb55YAQ9LBNae5OACMecm2Rx7Tf7mYafRwkRtcPAyGX3bLef3O+y+2fyLQ7QQsACiIR5/PI+F
XmAGBT6fAJOhaP0tNujd2G3MnNYDbZDcb97LtWo1ncUORsx5mmwP49igpGjo/qE4+XBpvyzI60Q5
AilIlHJhMKy33tCxgKL7Sokk8RPP4zjyWm+I+6JFr7Xy2AlMm67WQQ3lpBKn8bkUulnYKwkQlQRD
U/lngOjOI8CkCmPlYeN/ZoyST5P1Pj62wnUw6kPiHk1YqKH3pSkL6g0Vt8prBGTZWtknxcm64IS+
+v9LHL8HlH/ptgq6ZesK5HM7DyGvxIsYwSQOFlumDZ08Va/CKyH9J5V+EBA6n6pD+gcRGfcu9d47
WGyRb2/flgErpV1ulVJFHn19XnuzQoKbqhAs/PGNEaJUZ8I87D5MR+N1cohVvkQzBLAGqfF/5Rn4
l51KWzeXXorgjmlquKOwg67bMjMAuGHHOrXHri98Lx40Itpq3wdE5z96RaECrqMlCkCVjqPVgqEk
/ewXdcdPb0kwZ0YvJWm7uUk9Qcl6JnN7FT34xAc8YeOfz9EecWIT62in/Z7XcyoTIaJrJx4dJsih
jPgJrBx1nF+C9kkb7mjQWGjpRUBH/OKmXALdUPT2/qLacJY+1wahkH2b5/WObwPVdVKXa8nxVyNY
/AW0t0qycBbMjxE1UKQMpbvfL+Ojp0RusSj5o1z+susO0xR54qi4m7AbEsz4pGJhr1NEdJNY8pu4
/MtAdy8uL42zBdoPIc4Sr+EYcV9QRUEewUeUp+Sbjqfd6f16Cgn+NfJ/j8uz1SG7DDenqUKgS1k/
inPSZ9eTZW4QFau9msJil0G4iIL9jukab204eeBe7RHFRyPRDC3XN5L0s2q5RBd004IPbgp9MJYD
RFki65Hz7MfIJbiERObTe3Dcf5N1gD/NVz5P4DJvEsxstGryRmpn2r/28aLclGNlSNJdnqxqGVAb
zjaal93DaGyy0VfwSKraSqYo5nPUmd8bxKg/7mPpWE1TjIbdvEh1berdhRXxdK3ckpL4wFp8rRZb
wYdxoSWUJB53aZhDkqE791FK9TcfkDMTA5ugR0aVFbqkMh66B4S6ywFiUbrKQUxa+59RQvWlTOyk
actBGVJxZvWwo6EG1ZwNBDt3cA0w7JYVI4e8OPkwjA5dEKZ7agkTkE/bafkkC88xBxBc72Eskle1
lF8m6DOciIcNaTTKL0ZFyofs1+24fdbgfLnB6tMhXJsocFYVyitJBX0TvMc+2HU5MCCv58WmNi96
RgauuDvt9otVIIafeaemAcaD8HkWtbOkBtx+cDd/CE41RXfDDFoENYk+pcCqxhawG075EX2xpIh8
cBObkT6I/hlzZpT94g7sXfGmHa4Jw6SERAG0muTO6KvFnY3VO06tqoC4va2qxu9ugn7zrQZobRgt
pEcC8vLdMDCn7CiylAtKctZEBKhzrLhRWRl7UztV1C4riGjeL/D2F/y3gTFl5W1oSZXKai2mwF14
uxG7sTHsiGqe1Ac4/cpVOZEukGou3MAwE0lFTGwXkKJBSYVYtUkWONIbCQuZ4a0Hlo7NYajPjI0Y
WYqCo/iuqvPD3DkrZ//n5GVb8WKcKXCR7/VcZXeuecWECX9gNlidyD/8uVYhyHMW7vbAW5hjuAWL
PqUfKoCKWpbvkAEzgUc65enZZIG2DmcvatcOLlbxGlbcOZGZXphbp4yrv/2YI0t0Ly4dCX7Sunxx
EaXF5noOMqNIEvc5vYN4CJI0d9nWvM/44FS2jA9vsDYgT6yu/VIbhNODWVT4OjLPLT1wTzeAfRQa
T86BEfsXkWL2CWg2IRyOO7HvApga85IH+LQpIPTHOL8bdoSaMWAi1Pl743d+OI5INtLGQIBP5upL
pgKn8PI2odadyPqi9dxFXBpEKkPCvYPeReL2f5unQNAMsDIccav3nKNYk7xLEh7DWrk/aXdEB4BW
7Ct3az4678tIUg652jsP5i/xpNg+U1blj8Gg4zP3TRlKQ/VohKL1nZ+l7Jks9HtaSEzcGLKjPF9m
VwuifgNtraY8UhegOXpDd2D/VVv2ssxMiPbheAHZJIN4J3jfhkOd6L1UrQNn6EDb1G+sMRYY1zZR
aFbZOzimbtYQflzbOa26lz9ksO0Pf8Gkfrr5Ln4pxuA0kVD1xUWpYkcY63PfxWPVaHfsjewcoTmS
viViYkhMk1fmVkoRb/rR+KPgrfXH1rAex0b7FibDcsdj99b2u0/MjnoQ/mQ8Nsna2sAnZC9m6YLi
7lEzL7d0sbl14T4haHZ49bXWn7bvKeaXlu0q1cVJlSVTWEGliQ5VoW4f905KOD24kxjZuO4jOIWU
jupUvUp6cKVDXY4KLI93jWrsbuGxHENmSdslI2a1bsqa77NOpiFNO7Lh+csHlj53AlBsiRH0KvNd
BKtZ+SfKZFbXTMUAw+LThd64IsZ6SaFAnrFKmi9MhNP1p1U4jH5Y2qGU06EBznG1L5JO8AQDBM2A
JMuJ1rkHGI5uBJGU12+H9Bjdxmzj3++vIo//F1GM4UvO7kS8l0tiw+hyXfyGg7kOhUT73Jdsb77X
X7EJ7fLJq5jyrf9FIbujfJelbGtN0EEh+8plMYpoAkAhH+ba/9eXcKO30VaBJUBZ9BxfT8Y+/PzQ
6HexXiFPX7Qurr+hqp51uWu+iaPvtQvssiiuhechwUnD/VqbtXef4EbGR7w+akeOzBkEyVkoPhdb
rde3ZrXclMFwulpbcgr1Cm9uI+Cc8/blzFo4FaA2Uakq6xHHX2jbxBXD0Sg/7tDGuwBoix+VwRiT
kk9xTVCqubgKt73G3uBI4C3KTHZQWhhg6FRBhaDtXweiDf0hfaeV9g0jD460JUq3QR05/xCcaxSF
yYoDp3FpZh6RzOMCrJvCdhQp8OwWFGK4uDGOBkpJq+X9hZYwzV1+2szgNce9SFbmJfiGnK+8bOp2
5tiRihXa/1fpTnJWFuon7bGMr8IV03GgtW5waLL3q4JZ5sNYnVzYXCESH7sep2HYZ0x3+xZgq3Vy
BNn6LgUWIAeQ9hzXgazcA6ez8lPBw44lGiyHwBJNc4iKRyMpoFuDPiU+VMTs641INp9Gp67Or0UJ
PXNFFgjpdYSuzoOoTm/9kaBKL84vHkFa0IFjPLYpWONWVHTRCF8NOpsnm+037koHUmzkhk7dQ6r0
PLmF4yyoyOSE22BDFIIGByT+CSx0MGQbfAqlQN59+u3mOfIN9xyTXucOMjf9/VV1Nqv5Qjq/Hne6
SXjXk+G3kJvuSWu9b3exXSRkjOG7poGgJM3eQceQj2XxCY2UY4+y0mspJTSzFwFbYqlkk/9olaRB
sPP3732mYgxpZ4Rbv9JlEk5yPpOxsqxoG4FhdXIIvaxygmEux0vFrsxup1W5E+MyQ2HGw8z4ejdX
0tls+33yjnErzbFn+yTQJa76DjRghAtNztp+PN0ea4YG4FRHtVaUYmrnZQbnpMLaS0tsQN0fOC4d
BXrlB2Pdnb6TCCiBTbU0Fo7Qa0C907rbS4D7trZYW0ApIiI5g1JGOQVZifFdPzHb1QEC8vfH1auX
BaO12StYSfRa5r5Ds4RyoQJmPA4ruAgpzZfU1acflwfGQ9gle7gMhj9fQ5QHrVRWc8TtPkcuipNm
v8qaTfu0cwi0N/aQxUFdS5shueFs1KgbtGiqQSYW4aICtDLadWbvMMk5mzoIqoHrWUDjhVdctXWS
UFNRLfG5QESGAmKDi41vtd1gAJmNGn2sckcqeDFnwqxCqkEdsdf520PXEnLgmjqVdkH7RZwlNNVp
lurpmHdYL+l4p5IDd4Ek1NQbdQ5tzLvUZFTKhL7ZNJ2cUgEveKJ2prA24R00txfPvBMXesBc/HOB
oNwsTSnVG3y4euzh85jOCXImo+murpli/GWgevWn24Gj7anv/m+RoMGuKfd9RWEUzx3eQR7EFKtN
sEiYHpUL7D0fn1j6TlhdqlJjG1DHwXAFTJiTCtadrdvmuOaEpaFpVG0yAMQkWk4cIGk+pfcjpIBv
YFYO+gURd9r/a0bKsEnt0ul9DGTAv09e0geJDdS7+l81zsTbDviJZcmNpmWDIlPSuiadJ6pD7sv5
RG4ozuT5TdX2fonyAipmJyENgQH/irpWt4OZwVUywsq1z4o/zT0V0STZiWG867VKHDakG8kb8c9d
ksoQKGfYrXs5/I5M95FavNNdmD7weA9aoPS3PZhfmfYpxVf8Z/JaJLJZCl6gFyT7RLBnCh4EwQ3F
w3EyylSY/ENqy+zq5lgFGTE8WUKmbGtov1JopjgWC57E9eYtCXCc7WjzMEWWYRkhZAM38coJSsjv
3PE8zswvfhMSJ5VbFtV8k5PJX6IhbHRmXQL7MkHcsw89DKBMQEOBuHa+l7HTMRfSCuJvbGlPuMoO
oOpcSkp8WHG8n5U7b4YEACx7KHEbCytxpJWo0DaUIeZACBYhUpwEoNehcal2sqiMuqUsakAnebRQ
S8w+gUIVn4a0tQSwtx8z1ifjiPDxv3ZCpSNRAN4q/5jsDfE9r1RoCUub1/IGkwxvW7XKJ/MfePo0
J/oTXi+OxQOua+xvXNBTdbIMty2DRyZSd5QNS7bRH5C6P4LIvLie7Z9pARu0nHZYz50YLiuqz11Z
8ctwq0HvbmHhAWdAGjxB0KnkcUgnG2xp9Lbwr/dlJDGWBHOkWHQrD4aIMI0v/OmldB3zCck/Kg2S
qN7Eo3lZIPa51xLn2e3zxIBaYF35SzKqTemlP6768G377wcvoQY/yOYVZwA+R14Pq5l0+qwsgPod
FvqNbPiEm07LO8BC1kuunbsYfT5XRQk445SYcjLvcNz983FzXMWlAAe+Z41CTdMPVhMEpFWmRNdL
d55eebABPTXtBF092496LtfqNZN1AoAamasqPmWac/c9GlK62/0LVQ9XhORW/JA3dMmf4ReD6Dkd
S0AlGYWuUsiwj4Mcvy7ptKZs0Gd+dYpA2j0m8nC6ro06BQXaSgFb5ZH5xFbC6rNlDNi6jipFFtXh
eBb13C4q+Lwx6gKVgrT6XvOsm/2fAEk4IpKj0HkP0cA3X0lGecOvgYWUFhqE/ipM+xcr2tZ2cSfM
TIUxitFKncaKD4pzxfZVrRJOh30JL/0bmGiPyfx4WIl9FZGi/SOHgNUWQwgjGzzTJM70uAc2v0YX
LoT6NEPA+ZkSORcrcVNM+VqIb4sLSqxod8zY8e2+qNvfchoVVnWx7/XmTnDceUH2eir7+vvsNDmU
ZWJMC5HnV4AiCxaZ2oqXl0VLKbk43ZQdFaOgBQjogWCh519cyTdxOEBJjRa6+/+7432/ooBPIzSp
G09QKfhRQ4JnBi2y+8W1Hd++O1odLQNNGBmDWFI8dvZqdFqaBGZWNGm+WGzrqgDIb9XmdD1HT3dl
z4iMlq0/0RGwB6jpt0X8pKGoTzksvL5A1BnVLyVG/nceMZsnuRjoSG9MAzjA/dASSZMIlWOE8wm4
XvtCpD7+h2SCZz5nJr/JiQQKr8/JLs62J3xi89ySr32RqrEJ272j1eTLwrBKPs0ZJRbINhW2fSBL
xFlOiSopANH9KUGRVCeMFCJrV9J/QMoXjbl8LZ1CczAQ9kP2+pRcrllll7EdJCDiGJCHO4WdqeVY
DjEQ/W8rn8uC1dLryZ7gwTVef0nNhS244fGPlGBJZTRr0D7GI4enNF2Hiszh4yVYNY1GJy4yULtG
4fQN7CAzclQTysXimtKatBBCnAPbiBr7Q9VJo258oj09wMnYjTr7HuY29pnvN4Z5kLVFVOnRrqdd
mdxhh4AawZPxgzZAC6L0ptA0Wk0k1z8hQGYWjwQBPcc4sd2XB9vDWFI6CsEIoKwCPahDA4hJ1zVd
9phHrHTmMDt6sSpxXWYNGTRLXuxY2RrRWiAuSk3WJGNTp6G8uzE5aQmwN3HlO3fhB9ISpbh7O6Vd
YOFvgqre8x/IvrfBVCtCDXwW2TZ5++x6d3Qbl2tIECrkMMNpTRX4EgVxBqUlMZqKbaq+lNJuM/x5
uHvjJ6Fvg0UklQ/H45DtDN/2yZoHJqOxpvINMyVMMzmJZf8v5BkKrAqk2jU+UUX0DoSeFhFtapyo
oULDpJBoDxg2q3vHHFdzBFb8f6cE1CqeOo4ipn5wtjF6p72SilOxmBQa9o3UNQn2SZ8RpfJopcDk
IzgI6CMaVDrECLWmDQGKwsko08HQtp4v2HbIS8fQDogYKocEQot1PBNEFYPtlLwI36SNZrSXqoDi
BJbUt3+g2khldZL/mehRRvlNz8xwPMvBAU+PZ6V02Eg/kjLETxxcnCyeKmWC3iZeJQEMWAUh+6uo
sBf8VAz1MlWhCwytaQg/jo9gxlSbOp9pXiDHrIYSRXC+JEPaYBjkjAKcpmPYJVMr/Q+CbfbITv47
IXI00ctzRB+mQc3POnooNHo0G5qe/3WaDWZVXwlYJG6l8N+nLFEccma/wX+zDu6Mw32AAMtgapHK
CmxLcfKNSU01E1Ntt3ZzdU75rD1uJY8G4ynASqVkFFmyWsOr0DsqQW+tdwPksNMZJu3kXIHeTGjT
WVyKVC5mtfj5HTYDIpVJ9GwdUtSWmuD/PSP7zy4YziEhw3OrlbUxGKkKXXr17YW14UdlAhKnRxkt
Ye6vqkckRpxG42+SCEF7lbpy2nWwbcOuXrvC4EkLk59XsB7Ac2k5Xw7B6scwLkrJk3JOeM64op2l
+Rn+36emwLE50b0+EmSP5hpUbACoimvGSEqbq9/98FjhKzWte3xmFj2tubyrHd3Zgdh/maPNMT5F
4EBK/zYWIEVGkF8jjEAsHwLcHF6aYyWTd7he76CaqV9G6uJNwWGfWm8DXw3m6Xv1qnCWtoPA31zt
3W44axvmOzCnX4gUF3rGB2fDDqKNyBDNE/QYLlihHT3BxBwMTQkzVYLjYxelP4sP1mmXly7fPSRI
y24s+XWYe7x38LC+r9WuWlz8l7c3Cfz81xwr3En/ZOxM9fHf+VRbhTLRuvTk2CzRvlu9j6IbYCTM
SzFvziQ1F0oPpfLZkFwJMfzW8cWfyCnijfWBKeq0rnZgixIhBE3KlT9wGWdPVS3mNqtM699bnswK
1vaGd2+fQVL/gtjND2c3dJ4vX82Yc2xpF7fpsmbLqoZkK65CrKAGGnQFK4oHyRkoOPfDK+HWOgPP
0aJFKE7HAfVDfjaIau30daLv7/mEg+7LXPsGLXoxG5YNeYD0S+DVu4HzJNuIbb/WRp6LzMXXSJ95
lofst1ACplyc44o76XXOJniPIQhQEJamTYfbeOUcEjUFc4GnJjjtZ/Rv/0hTel+C9FWfGu0D1wBN
nGNI5gN1wO30vjnRNYGZq4DVqtQ65EPTaooF+r7bf6OH+cvis29owFoIwCxxUGyvfPLqGhh9rjpd
abiRLMGUbesBY3WYiKsZYj3u7PVex2NMDxb6Xv0AkC7YpKsIjSZrQwX0FgmplscpTH9gkH2Wi/6s
JVIo3CaKp7Eqg2EP0xsM6XAlROKx04H/glJnQbm7vNmRvbWtK8avpwp48PhBbdOYY7Kzz+RyZmHZ
T45cdo4/ytAswaiOY3G+mGWxvZ0JdVJXU0SzTJtAjOaLeFx81ZpXysRMViufGPmgIqOaZEgdkJlc
OibKSUFIzu0vcPooVgWYMEk8+e1O4/fDqaBOW5g5NJv8vIpanc1ReV/WbWco78RZ41WyYBStZu6y
T9MeiRt12Zh7MW/cCiVQ8kbL54TXnze73s+3NN2JQYKZpZccX6iWQDQqCiDILotSN4zX1uuyZIer
tgYUS9g2SxT35seGuRWktD18DyYjgGiLDVf1Cntkw+ic2zUfCOGy9dcenaAfO36mrdhJS6vq205h
k6Ldqa/3YMXOC77bd19SNuami3l2FhLWyqNNEyUpiAgw3lLE7q0UA62m8CAafa8n+XP0uW2a3CIm
M/B+Zp363dKue++gDRO4lD0DYvXUXw3D2jIoO6frQ1HX2J04zJ0ctf2H13uGhd1neW8pY06xZmhs
iq133/XwomxWika0BZmag2OlQqRULIzBTL0hEZR8YUDE63IjL78dqyy767MQrhcN05Wlzi/cnUyi
7u/tJKQP/FTbIv/kLTegX27fWSfQfEhEbzyrXKfn8CXvI5NXVsSv24me87rXUnGR//yAT0OU3X8k
oCexEJIoLj234RKNCGgxz6lUULDdr0r+S5J98GQmOCFrdGBL6T3O23mSTQni8r54NJDGyj54T7M3
A60HjxeSSla22HZw+WqpsfkkTecOWQ68+7tt3zJiHHDREIEDMc4r8mRSy6fzWIF8pPywxmyl1Iyq
/Gm/+jB9D0FRrJun2vgiHiaijEebCe/JqQ6Oc+78ufQlvV6bQB7B+0oRw/62xLMtUX0vqB2tNnPw
+9iDMnfjRFjbydq588WV+0O2QN0WGig7Ohs/8uEqLciYyronjKw9c08JfAsiwXynF+1P/Mzdnapt
fg4vfC5Yq8TjdMW/0qIcVNRv/Nv01STegh5Rgiq5lKr0FBg9oixskjzVGDUfUXuNCL1m7gzp6UlH
Yi/9S3sUkOfAwlsMdSgTlekW6kg6rcRwx2PAp4mEwK1fLnUaLvLG3R7jxa6+DJuPCFxxjq5tcaYz
RTiYYHEP+wJW+Zw1DdaEZR6o3Y1VBiUH/RtQ6n816j2ot1up64mQUgIWschJTNhFW68Wg5mfz+zO
5hwHxsJw0V/NFSZng9YowgKbY1HiTW70GVwAAvJrX8TiueBIoGffzXw0haXZs2EBJlbHnUBnjmQx
0s7U7fGEkf+/4wFVZwSq/bpWpdxoPzOVrkOKpXYKPB5nB/vuAl7C5PBTHmeGCUaB6MrZV9zo6oBx
zG5O3CUWhORxutOaAAFFPBzTUTun16enkDEJW1/YNTn/t6106uF6CxcyBxiGLI6cZbxM9SRnfuc1
Uw3BcwfHCpUOC+7dzdS467dGVrmTzeyuCO+rZ4Ivd6oidHQ7xZ4v
`protect end_protected
