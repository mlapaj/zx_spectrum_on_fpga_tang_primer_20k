--Copyright (C)2014-2023 Gowin Semiconductor Corporation.
--All rights reserved.
--File Title: IP file
--GOWIN Version: V1.9.9 Beta-4 Education
--Part Number: GW2A-LV18PG256C8/I7
--Device: GW2A-18
--Device Version: C
--Created Time: Fri Dec 29 22:53:35 2023

library IEEE;
use IEEE.std_logic_1164.all;

entity Gowin_pROM is
    port (
        dout: out std_logic_vector(7 downto 0);
        clk: in std_logic;
        oce: in std_logic;
        ce: in std_logic;
        reset: in std_logic;
        ad: in std_logic_vector(13 downto 0)
    );
end Gowin_pROM;

architecture Behavioral of Gowin_pROM is

    signal prom_inst_0_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_1_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_2_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_3_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_4_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_5_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_6_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_7_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_0_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_1_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_2_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_3_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_4_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_5_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_6_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_7_DO_o: std_logic_vector(31 downto 0);

    --component declaration
    component pROM
        generic (
            READ_MODE: in bit :='0';
            BIT_WIDTH: in integer := 9;
            RESET_MODE: in string := "SYNC";
            INIT_RAM_00: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_01: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_02: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_03: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_04: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_05: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_06: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_07: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_08: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_09: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_10: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_11: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_12: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_13: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_14: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_15: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_16: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_17: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_18: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_19: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_20: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_21: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_22: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_23: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_24: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_25: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_26: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_27: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_28: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_29: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_30: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_31: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_32: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_33: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_34: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_35: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_36: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_37: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_38: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_39: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
        );
        port (
            DO: out std_logic_vector(31 downto 0);
            CLK: in std_logic;
            OCE: in std_logic;
            CE: in std_logic;
            RESET: in std_logic;
            AD: in std_logic_vector(13 downto 0)
        );
    end component;

begin
    dout(0) <= prom_inst_0_DO_o(0);
    prom_inst_0_dout_w(30 downto 0) <= prom_inst_0_DO_o(31 downto 1) ;
    dout(1) <= prom_inst_1_DO_o(0);
    prom_inst_1_dout_w(30 downto 0) <= prom_inst_1_DO_o(31 downto 1) ;
    dout(2) <= prom_inst_2_DO_o(0);
    prom_inst_2_dout_w(30 downto 0) <= prom_inst_2_DO_o(31 downto 1) ;
    dout(3) <= prom_inst_3_DO_o(0);
    prom_inst_3_dout_w(30 downto 0) <= prom_inst_3_DO_o(31 downto 1) ;
    dout(4) <= prom_inst_4_DO_o(0);
    prom_inst_4_dout_w(30 downto 0) <= prom_inst_4_DO_o(31 downto 1) ;
    dout(5) <= prom_inst_5_DO_o(0);
    prom_inst_5_dout_w(30 downto 0) <= prom_inst_5_DO_o(31 downto 1) ;
    dout(6) <= prom_inst_6_DO_o(0);
    prom_inst_6_dout_w(30 downto 0) <= prom_inst_6_DO_o(31 downto 1) ;
    dout(7) <= prom_inst_7_DO_o(0);
    prom_inst_7_dout_w(30 downto 0) <= prom_inst_7_DO_o(31 downto 1) ;

    prom_inst_0: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"4845BD5B243DAED2B2489B313A35C50252AFD0FFB76FEF342335FFF132FD92FF",
            INIT_RAM_01 => X"5372B72B484E2F2664B735B69A5AB532B086BA4C62AD6D56EECBDB6984B25145",
            INIT_RAM_02 => X"DD6E630C15271E48CA801988654FB501D5393392EE765C1EC95C1E4D86F18A96",
            INIT_RAM_03 => X"17F7F5724D40707E6FF30002982023020449B4680C45D1CFAD8EB30A061DB8FE",
            INIT_RAM_04 => X"BD52921D249E377EDBD14EA309EEDAA57DA85F55DBB7048A69A4C801013948B6",
            INIT_RAM_05 => X"5E2B1A3E16869E1D37BCE906B82F401CBD467617DB34D9E0C80B5E6E10063EC4",
            INIT_RAM_06 => X"BA611013110188547995B108BB2DAE76F4A3A0D98845F9248BDFA45E10CA403A",
            INIT_RAM_07 => X"D0734B461A36980411EB2A6C1BE76029258777EF227A8F6E84F74C4436098F67",
            INIT_RAM_08 => X"60A229B98541E6FE734DE2280A9B57FCD5A9BEFEF7CDA5ABEB44FD73D2794D56",
            INIT_RAM_09 => X"84735325ACC969B2EAE10A1478D866FA67DDEF7BBF75E6958B6D02DC6D0F8076",
            INIT_RAM_0A => X"7833830C7B2C7AFB8A8D203C312306DA0E72641FFB93D79B5EC04F44AD55F4B8",
            INIT_RAM_0B => X"1C387A7970C7F3E688673CF5975EE3E5FF105CFCCFAB725D698FB088B063063C",
            INIT_RAM_0C => X"96CE81973CB55590446D599375501366EC343561BCF83357F8823671393B278C",
            INIT_RAM_0D => X"8CEBCB187AE5D44ECA689C9BD4E5AE544DEA7E90D186B9F335F3223877AAD541",
            INIT_RAM_0E => X"BCCF19EEF299751C919C9C13C6FB9ED711AC4DA7D947CC79E9B6323EF6CE6263",
            INIT_RAM_0F => X"763DD7AAFEED3F4AD4EA7491ADE6F14E6DBADD0F090A8DF34D7BAD35DD2275F0",
            INIT_RAM_10 => X"37309C08305A10187707E3D57DDE4931F1D9E97A8F378981ABBF8D7B6B7549C3",
            INIT_RAM_11 => X"9467DA6C480E6D19CEEA8451CEFA88FD70E7925B0302F877F87FA833FBD147E9",
            INIT_RAM_12 => X"99716B8CBAE953D061FAC3D6337D5BA4D6D7090929944AB6FA3357801066B658",
            INIT_RAM_13 => X"F331598B364EF27516CC49A4662C5E5C92ED140D9637367A7833AE4346982375",
            INIT_RAM_14 => X"A5875745B625C6CA7A7292332492D139728A689DA1AE78B6B44CE4F4A4EA5A22",
            INIT_RAM_15 => X"CD2E1AF14C30545297A91BED3AEAEFF8F696B5F4FC80BC6B1A2559492E9198E4",
            INIT_RAM_16 => X"75B74FB9AF7C1A492952F7EEAA0E7CF9FBEDD0FB47EEFDCC3734B816F355C913",
            INIT_RAM_17 => X"88537A811D4EF6CD9668CCD3E2E7A8041788DCA5F7E08AF52AF527607BF06DEB",
            INIT_RAM_18 => X"66591A35ADD26B6B7E33CA56E9A4759EFA7E68F98AE7CE9507755C74C430286A",
            INIT_RAM_19 => X"56F9FDFE7D64C1F4E1F5641845CD17E836B97780400C702723FA8E7C7BBD6F06",
            INIT_RAM_1A => X"0A01FDC7FE2CBF038A61DEA5FCE2C10C8F35FBF80C05ABFF4B6935287B125E8D",
            INIT_RAM_1B => X"605D53A5C955D5D1412F8361617A54446971FD187442A60FB04457857BECC312",
            INIT_RAM_1C => X"CE4B65409D6F079D709A56C38DC3BCEF07459A416EB4E8F3D73CC714F4333AFE",
            INIT_RAM_1D => X"04B57D8E0D755851232838F9B5348838530D7AF95411555D263B8CA86A5D29D7",
            INIT_RAM_1E => X"DF7D7BF31C6072BFA7993996AB7DD2F3EE4009844CC9D6CF9E583AEC48A52F29",
            INIT_RAM_1F => X"1EEA3633EFEA856D05BA968C1B3C30CA1788DD95D16B8F914DDDFC3EE5C69945",
            INIT_RAM_20 => X"95DE707778B17C2379847A23AE6B8BB01F36F3F44A8162566D9FB15DE7CC83F7",
            INIT_RAM_21 => X"EEC890579E95D5A0A546CCCDD48577558ABE7CA36EF67A70F6A8758BDA052D5B",
            INIT_RAM_22 => X"6BAD12FDFB527EF4F87F4A23EC13CBC0262D8899A3A290F04F41C1324045B9FC",
            INIT_RAM_23 => X"85287860729C77B6C68CAEA3033A6E84D67249B594C407B39C68B4C1C97FDEFC",
            INIT_RAM_24 => X"CB76FAB179E9619BC7E7E9C9FD801CF87DBA1EA496E829D4E62861E1AF436A75",
            INIT_RAM_25 => X"65F627A15E1057ADEE7B9E27122A58FF2B98B1EA560390C7E8F715861814E04D",
            INIT_RAM_26 => X"0004406BD60A023AB063D4E5966EA41AA997F5A49BFCB0657A9732D28EB8217E",
            INIT_RAM_27 => X"4ED4AE2B1650D21EAFE01E7099EFCA3094FD4D705CF6B84AE21583E13385F865",
            INIT_RAM_28 => X"5725EA43CE18F187A1DE4DAABEA97963E3A7A96B8B7CBC095BEB7CE46274D9AF",
            INIT_RAM_29 => X"3C563C8B02C8CC39C64DDCEA1BEEB5E7353F93786145598FE634EF1000179B34",
            INIT_RAM_2A => X"735AF87DAE59FABBD7DEAF8717F2B72F428F5E37E5D6E13157B99CBD2D73B9C7",
            INIT_RAM_2B => X"9555AFBBD3AEBFCABFBBED7A5C5FE9BD0E6A91C6E7610042695EEB08D8881B1D",
            INIT_RAM_2C => X"C5595549AC64787878F5CE14C664CF9EB0CDAFFBABEF1E83358371B9ED96E506",
            INIT_RAM_2D => X"CAE30B9FE6AA29FFF6F72DA73DFE4F7ACD39687B9E69C5359E9B991F0746EFFB",
            INIT_RAM_2E => X"EFEF92C2FA4D8D4E4AC86C277338FA37BCDD9D47781EDBAF7FC03C1BCD23D0AF",
            INIT_RAM_2F => X"E629BDF93D7F5B5BAF92FBAB477E9B315DB5A310CFACC7408DF9A544B1E57AF6",
            INIT_RAM_30 => X"3F1BF746FBFFC353E37263FF38A796EF39E3FD7DFEBA7FFEFFBF17ABAF09E909",
            INIT_RAM_31 => X"636CDEB4BDFCAEEFC61DFFEFB7E26262DEF2CB9F71565824FEBF3F7BDDEABB59",
            INIT_RAM_32 => X"FF9FFF6E3881C81AFDCF2257FD4F8ED5257D0E9B800726B646C8A8E5012F76DF",
            INIT_RAM_33 => X"4E93FD3C1238FFAFBD7FDF567FA8FEF024F33AFD3AABC6B105EA80272D64895F",
            INIT_RAM_34 => X"47B2AFF5B87AA26AFFDD317DEDCFBDFFE1A0CAD3B58877DD2F647F7DF748E7CF",
            INIT_RAM_35 => X"6F6DFFF29CB70FFD25A59DFFFED7B3F7E8B4CE6FFF3EF9CEC6BAE57ABFFFCEE6",
            INIT_RAM_36 => X"AEC4837C2A5FECBB94C1C969FFDDFF79BFFAAFDCA8D748399ABF75558ADD02F5",
            INIT_RAM_37 => X"DDE6FC8EBE3F9F3C3DFC6E8F07BFD31D50660B1E0B2506A533CE0E340C7C745C",
            INIT_RAM_38 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEB9A44CE0EEDBBBD391D3128AAA3",
            INIT_RAM_39 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_3A => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_3B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3E => X"8000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3F => X"3C00000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => prom_inst_0_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_1: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"AD5751BD429B4F61318427560CE39D492990013FD212181064E2FFF009FB997B",
            INIT_RAM_01 => X"8C6AC955A8A6140421573E413CF5A80AA1436D8B4C31A2AB26D2A61CE834248B",
            INIT_RAM_02 => X"6CDEE7468681D6C31E4991CA3736E9ACB7531EC6D8BBCD453718101EA25D7927",
            INIT_RAM_03 => X"15408676F600F490FAA59B488C7998CC8CCC28922AC62644EEBB432EEECB51B1",
            INIT_RAM_04 => X"DDBB7B207EFA17098E07684801BD45625A36BB62220506E171891964A31BED22",
            INIT_RAM_05 => X"FA4F91915C6AC9D8570C292F10848189906127BCBE06FFE92DAFB4AAFB240D88",
            INIT_RAM_06 => X"4CA272352720BCD900A6D79BFD9D0595EC0D044ABC8CC28E9AE946E3D2000A4E",
            INIT_RAM_07 => X"9C8CA06AA05B63C89A59A3E4E80807B27A70B0006624C4AC4A0995CCD8CA2082",
            INIT_RAM_08 => X"06C78011F78D8B82E59F0CD4B32D6801669BE3EB0B96960DFF152005EC7C16CB",
            INIT_RAM_09 => X"3AE624C94932927924D20024CD638A01C8620023319662D80E05805625BC4A40",
            INIT_RAM_0A => X"8366123AA809AB30B47977571C5D70397A93C723106D0A2C254714359DC7C9E1",
            INIT_RAM_0B => X"39BCEF6BF4D23532957455F1C80115524179D59C4C4534DF7296991146CE2450",
            INIT_RAM_0C => X"9E2DBCBF62498A769883D7218899245CD18AE49F0146517422EE475D520029ED",
            INIT_RAM_0D => X"E9969472A81B83113144528F831AA6C3221E137C1E9C670E26808A894013828D",
            INIT_RAM_0E => X"9FE2D1F27443253D58403577C801AE23371F00290A17E1C4A40258BFD204230E",
            INIT_RAM_0F => X"20721F982534A8179F13E2C6328CDE7D2A73087D3A9314419022103DFF767776",
            INIT_RAM_10 => X"7DE6C2ED45D76325CA2A8E198859334553AB02945CAB1F17C142288008073004",
            INIT_RAM_11 => X"0644C9567C0BF9911B870B989C59330089AA4C8065AB1B11132213EE0FD83081",
            INIT_RAM_12 => X"6AA394A8644494895569192AE42AB508290A2CA59B4D6EF213548EED8642F231",
            INIT_RAM_13 => X"71163594CEC5863F0F56625E221D6B8180848C6B2BE24AA2AEEE5D187201CAAE",
            INIT_RAM_14 => X"198817644F293AC1946061117122A39D8841818C1389D51BDAC5491819025165",
            INIT_RAM_15 => X"27929938B8E10530250877A4998D0DF0004852125C20CA8D4279881E41208B14",
            INIT_RAM_16 => X"5E1384C93920A16C9B696272DE7A2948BE8AFE81310146B8AAE5E549FA27EFBE",
            INIT_RAM_17 => X"376E511217E00B624A46BA2E4CC10B729C326F710F24CFE78C5E63F3034737CC",
            INIT_RAM_18 => X"EFD5995634050D4CFEC166B032BEED5553AF0358304080D9DD0A2E9948593830",
            INIT_RAM_19 => X"C80CEC08A7F5F85CE65326632B4C4F3920019A35AE2AEB3A1131046EE45B81D4",
            INIT_RAM_1A => X"5939FC47C933E1B0AEF12AC84454CA47B00A6BEC5402AA08B5106E3065602454",
            INIT_RAM_1B => X"EF30312A73337CBAD4838F42A3293859CD169240D8E652F6D72D8D19D56DD767",
            INIT_RAM_1C => X"E2E0440C6CBD60741FC178643A852D4A2A0627C688D905B882524E191E7951EA",
            INIT_RAM_1D => X"36E0548D65FF9125A765F0220F6EB9D1B318244CC6CA2CBC9CEC6979C14EB28D",
            INIT_RAM_1E => X"082C891C76A4845096304A0D8502080C1198921998821D11C29CA830C3374992",
            INIT_RAM_1F => X"35C65240B61076066A23CE4CFC5E76063A1C2AE07DF555007338BDC080EA0C23",
            INIT_RAM_20 => X"639303AE5376F664C7125632C19440CECD5740C77849D937472B202579964F60",
            INIT_RAM_21 => X"14E5DCCAFE50CC13922A5B149C598A621F80C24D215291228844E7F33F9763C6",
            INIT_RAM_22 => X"21D9DC46629BB376E97F2C7BF8C3A218EE79DDBCF886B2BBDE702F71B38AEC69",
            INIT_RAM_23 => X"6EE48A1CA6430860DE613153615CAF4C8D191004CE9C6105D8C6795B6484467D",
            INIT_RAM_24 => X"9F0120108829220B230F44550832C1022530CC13C4C30D8254ECA5200A194126",
            INIT_RAM_25 => X"C0BED5FBD379F904A41BAFB6BE4EE9F6E8058229DD0C354F03CA6C4D8B6C16A2",
            INIT_RAM_26 => X"5621E625522D34519BF2C353F8AA030B9109C2F9686AD3AF57AF3016D9160354",
            INIT_RAM_27 => X"5FFE6AD3343986C4103935236B6E6E11B940EF46A8FC06E6872A6929D50DCDB7",
            INIT_RAM_28 => X"7740114D6B08228BCC693FB12CECCCD2461586069445ACFC910B1241434622B6",
            INIT_RAM_29 => X"C08C4847914664518E27EF7EB9C870A226AFC35BEDB651840466400D4B3C0F87",
            INIT_RAM_2A => X"A807C3A1110211AFCA2A142F0BA928156D142250438143D339E4E2079F298493",
            INIT_RAM_2B => X"7FF29C990C9E66273CC78041192D03081CC62A8A0D8CB4D9CF2F2558131A78B8",
            INIT_RAM_2C => X"527CCD419525AD29AB7D372C0B56AA0A065F8BDC905346478059EC8280192068",
            INIT_RAM_2D => X"12D552A8A0496EFE3AAC6F34739A94E798101823148D811212E9A349CB219049",
            INIT_RAM_2E => X"01DEC1A54696B9912E8B0705C8587D4F7D36C863897BD3102AA663B819B55B7A",
            INIT_RAM_2F => X"2C05EF54A3C0F7F5F017E03F5800377CCF6E493C84E8F56441831087370A0848",
            INIT_RAM_30 => X"100E0A7211342DF02958046899EEBE6E491299A09312778193FF3D7FFABA8000",
            INIT_RAM_31 => X"1A94A248414CE030020F207BF040A06A3DF993DEA3823423F405294A52014565",
            INIT_RAM_32 => X"AA0AAA22B1C70003F542A66FD1F1CF9D4578315F8C1C6FEC4FEDBDF22CB20482",
            INIT_RAM_33 => X"00D988737BBB44C414210118C673B0C1BDF76C499226F78FF41A0AF7AFD3308A",
            INIT_RAM_34 => X"6087F8B130F04418C0A1C082FC005843F5B42CADD9455ADBD328C13219110DE1",
            INIT_RAM_35 => X"54E09A38775020189010680840800297C31282442326D008D1F2351A89FFD7C1",
            INIT_RAM_36 => X"A0D8E36A84D5C61285128845215F8F8821C308E368283D8E2B42989C04A8B513",
            INIT_RAM_37 => X"81F3167814687CBD683E54D44555E6C95B5F2A72C0C193C6110C0221A448D0C9",
            INIT_RAM_38 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC4503442C4F91309238ECB252072",
            INIT_RAM_39 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_3A => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_3B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_3D => X"0400280000003C3406303220344C403C04001000101000000050627424000000",
            INIT_RAM_3E => X"80000000424202423E1E3E02304C3C0C3C7E7E40403E427E3402421824347C1C",
            INIT_RAM_3F => X"4200000042000000000000000000800000000000000000000000000000300044"
        )
        port map (
            DO => prom_inst_1_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_2: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"9E28CC30C7C2553DED3378D655AD194B2E6C1CFFED700F6713D9F8F33EFC361A",
            INIT_RAM_01 => X"71A553CCDD8ABA79BD27B7AF735ED2D34F1EF3A81A160C9ECB1B1FAE6EDEEFF9",
            INIT_RAM_02 => X"F6369572C3BB8AA1984A8D12F776E224ECEEB21F97FCD6C0CF17A044EC2BBF05",
            INIT_RAM_03 => X"E51D405CAF70F622DD4599602D7910DCAC8214B2A4202510C593202C8B164C8D",
            INIT_RAM_04 => X"34ABEB9DFAA4853910C9965C158947081CA41402E8E65478737F73BB629AAE2E",
            INIT_RAM_05 => X"F84DBBB9878C55457324E92D3DAE91D729AC76BBAD4C6EECA74DAB5EE9A175EE",
            INIT_RAM_06 => X"D7779D7B79D1C75DF87378E98719C1AF38B1B801C71D180CE86370AE9C2BF38C",
            INIT_RAM_07 => X"973FED2E9BEDBA474B70B121A8D60F3B4EE3F1A238FB3B730EDAEE74EC632DB4",
            INIT_RAM_08 => X"27271C28420E47B8DEC74738FC3EDF9FBD40EC09FC7B4D3A1475BE433705FB5F",
            INIT_RAM_09 => X"3091900604017933442359491FBAB63F346F0C5EC8E3A531984B09E605A30A06",
            INIT_RAM_0A => X"5699692496359B8E67A7E74D9A0FC504C8465638CF74A1AF9185921A7D262989",
            INIT_RAM_0B => X"352CD1DAFC910CC504334DF9E6F1F4F30161A36293CC5CCF1CA13994ED29D34A",
            INIT_RAM_0C => X"F00030AFDB7F22E68CBAA4D9BE7633D3B53E90E4B124422A2A4454BACA5A8DC9",
            INIT_RAM_0D => X"D195D748900C29DF7F381280A9738CDC3BF5BBF937D3A4D99CE2ACCD97CEF2C7",
            INIT_RAM_0E => X"F1A8CCFC0C7A15BD9E7C2557CB00BF2584E16AAD13D7EDB525A85ABF90C0136D",
            INIT_RAM_0F => X"386BA04EF97A3F8551DAD9D24A8D259A03ECFF5AB81B1C31DFDAE10100544F8C",
            INIT_RAM_10 => X"7D94E6ED80D6722F3989B91E31C63B64C363DCE71A861C14382E270FC02878C7",
            INIT_RAM_11 => X"293A130C900FBA4EA70D2BA25B343C5B026D8E8766A4E4267CDAEC99E830D230",
            INIT_RAM_12 => X"3B9DDFE4F83A56E124BF5BCE9B34FCAA67E49B3A42E19184B6C9F07349210436",
            INIT_RAM_13 => X"B755D1CBF0DCF6FD40BEEC16EAB4A6D16839C98CBE9DBB42FC69FB709F8E7999",
            INIT_RAM_14 => X"5ADFAF6726384795A7656B753D2369B9EB5595BAA722012DF8DCFBF15BF46D6E",
            INIT_RAM_15 => X"3AC884B1E69101135CD080022451F20884CCB9CD203C141402A5AD293C3BABA9",
            INIT_RAM_16 => X"0AD005E832924E92429C091D167806C10041AF32DDE13A669990457D098CC2FE",
            INIT_RAM_17 => X"9A2921ED6AA0CC8387B267B9E7A182720833CEE061E6450C8E4A72E3C087F21A",
            INIT_RAM_18 => X"89A4D43867379AB880C1ACE279E8DA4B3A9063A0B320F65E536B8EAF9CBB9C76",
            INIT_RAM_19 => X"20C76D6362915156A7671331CE657011862E594E46A6D99992E2D640D7668693",
            INIT_RAM_1A => X"3AB1F9007B8A7F2936D16234F9BF9B6BABD48FCE74047C1E738C5B303E815BA7",
            INIT_RAM_1B => X"027170C5DBCC2B6AD72B8E4CCC94DAA139D8BA64E3384337426E7F274CC88A37",
            INIT_RAM_1C => X"144A4566F47B73C95BE6CDB9E664D536762E9224D70F9A5C374B4D1CAB8DF527",
            INIT_RAM_1D => X"7DA5F4A8458A9451315B681ADA9AB0D63218DFB77D3353C32837E954604B9D98",
            INIT_RAM_1E => X"F7D3C6CC8C7841AB49CC538E8A72F2E73C64D2DF3662B19407D7D299CBEDEF3E",
            INIT_RAM_1F => X"77A47C739FF6A22B8B5CDC49E748E9C739BDE6756DB4D22437E74183E12400CB",
            INIT_RAM_20 => X"177AF49DF118FE47ACE3344964FD4ADCFBB543F7729CCB340866D1157B6CCDDB",
            INIT_RAM_21 => X"D6E60DC661155EC9E80F8CEE659F19CC554B2C67C33EDCDA63BAD91B7D1842A7",
            INIT_RAM_22 => X"00FDF3B9B8DE5B76E97F8D32F0F39E4CAC68D9BBB68EA3915F6225F932CAAFDA",
            INIT_RAM_23 => X"441A0CC068A0823F8668A00621B779DE35FEC004050469F34866AEE766743D8C",
            INIT_RAM_24 => X"DA00FADB1D3A630BA18050635DE7DCB13B9B86E0CE6E08DC46331A352F716E3C",
            INIT_RAM_25 => X"A5D31B86A0288D29CE2EAAFF86A6A9F3000082293E6BB54F06698ECCB199973E",
            INIT_RAM_26 => X"D972662C0D31E34E63B31CFC6EB4B35A69B67D85489E62EA99899A94F6800FDB",
            INIT_RAM_27 => X"7FC8531A7A319F3EBFC1383FFCDB0E09BD288288B078B4AD220B6FA934CF6187",
            INIT_RAM_28 => X"96450B74E95A860FF3E434C65F1308F16F92395816B914F0CE870C1323347A4E",
            INIT_RAM_29 => X"7D8C4C59396600DC0C420495A0D987501490002BAD38012E20620D556A230B17",
            INIT_RAM_2A => X"315502751655F60070E6B2C50609369611365AD1E3352327320331A51818030C",
            INIT_RAM_2B => X"AAAC4802B74190FB007C0C0206186AFC1B3A2A46864F26118ED1D03ACB1062B7",
            INIT_RAM_2C => X"E73D9D6D2C265859DB844C2C1952AD10241100174FE0444E6707D80A098D8585",
            INIT_RAM_2D => X"8CF14A288EAE3BFE00FB2DB45080D4A50C58263A3B398DD51AB9CB554ECAA7B2",
            INIT_RAM_2E => X"03AD0025F0D509F63202D877ECD8BF8005451F7BD37367CF0BD9B79850A7D80A",
            INIT_RAM_2F => X"6C60009CA281AEACDC1762945981B869F93D683EAF4AC7EE52412E85B60B91CD",
            INIT_RAM_30 => X"2A191E00538FC8A5004036A959ACB7A463D23E419EA06B744006385455A71250",
            INIT_RAM_31 => X"464C92242004E0AE8518E001D124A7628010115D23C30462FC00A014A1213358",
            INIT_RAM_32 => X"55B555C2278100000A24804D7D98EB98602733818A12094F0B6515022CB40002",
            INIT_RAM_33 => X"4683814663FB910969D1D631A952B381B7F635A33FD38D5CF15DF47D057F7FF5",
            INIT_RAM_34 => X"6A855EC94CFEC4E0172C59A7D054F8F9F4356C312C204E40B05E2059407C8DC8",
            INIT_RAM_35 => X"B38F54EB9091AE3320201EE395AD63902282A031CE3E87CC902954AA515D5D6B",
            INIT_RAM_36 => X"2E5172E82E845070000A846100500E84EA1803B8B07B99E1DC75BE6419674597",
            INIT_RAM_37 => X"A111466C9493A2A7CA2204102414CC798BF0EEC2995A4814580BD07585585ED9",
            INIT_RAM_38 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC25019C244097049C2B2DC8D93C4",
            INIT_RAM_39 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_3A => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_3B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_3D => X"0A1028440000524A0A4A4A204A5240460800100010540042002064547E060000",
            INIT_RAM_3E => X"8008004042460424402040024A3242124220044022404208520A4A24424A125A",
            INIT_RAM_3F => X"8102080042447C443C0C3C402004FC1838787840407A00707C02487E44487842"
        )
        port map (
            DO => prom_inst_2_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_3: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"CC8070206B8245AC240020752EBC2BEF3E748D3F8F360C239C4AFAE93FF8775A",
            INIT_RAM_01 => X"00812F408CC6501331852531B04480021D9220D4903A41404312032840153FE9",
            INIT_RAM_02 => X"B383E6E7C3B310E1F7FF595C5DF6F0E9A9FFFBE16D3FFBE82C1E0051F1E060D5",
            INIT_RAM_03 => X"C1FFFB3487617BE24FD79501DE05F1A341B89EC82FD5702597FD866639C0DE08",
            INIT_RAM_04 => X"47A8EA413A2DCF0BFA8EEC2318DBF3C4711871B3BC0404EC45252A485234A663",
            INIT_RAM_05 => X"1D2FCA8DCB43C5356BAE638588C302868CE1161CACADFEF7696F8C3AA82EC16F",
            INIT_RAM_06 => X"FF4DEBFBDEB376DF68D5EEDB5EB4D5AB5B39745D76CD8ADC59CB30C8AA33E155",
            INIT_RAM_07 => X"06ABC52D5DBEF57EEB3311A9D85D253B44E250E1566BED57C6DFEB2ABFD1ADF6",
            INIT_RAM_08 => X"D7D77EF5E2C6D7220BE64B3C6E9EF22AFDFCC8005C2FFFFA3AB9AD1ADFC0AFE7",
            INIT_RAM_09 => X"DCD4560015805B13AC0290001EF826137E4EB867C828D9777FFF47B6903008DD",
            INIT_RAM_0A => X"1C9DCD8EBB9D36AF570CF25CDD16F645D1DE9F9EE575E2A2B91D5659FC131CE3",
            INIT_RAM_0B => X"CF133BF47B9D3DA46DD6DBF3A8ADCDD3DF1176D2FE23447DFC65E1DD7BF3BE5E",
            INIT_RAM_0C => X"F0A09C47F23F20FE2ACFF5FD3ABE6167E5FD36E1D9735BBD5375C1F79BD0424E",
            INIT_RAM_0D => X"3497229CB9044B6E7A7861A04A712AAF29EFBD393727F1F3FC2AB1E6CF571457",
            INIT_RAM_0E => X"A8BCDC266655185CC45008B39EFD1FA6E9F5E816114F93E1E7A2A27C72C7349F",
            INIT_RAM_0F => X"FD5CB07B6C729B510A78BEC5F7C7A1E7809F1976D0DD3615C1D27D2DF596BFE7",
            INIT_RAM_10 => X"63B065F7D671322D6BFB2B8759433929CEC27E3FD7741292A4A5AF02703CF4E3",
            INIT_RAM_11 => X"DDB3A42AC80797FDEF4DE3EEF7ED8C7307E4CE6A6317F7BF25D077BBF03AEA33",
            INIT_RAM_12 => X"59BD7F8DE9FBF27A65DE5245BEBC7DAA0A70DB7240B0D136169D77D649A39EB4",
            INIT_RAM_13 => X"21A40982C046D22C10146484345CAF7BC828BFE79DFBE3C4B1CBF660C487EBB7",
            INIT_RAM_14 => X"CCCA0665222D038CC873351A21B23939A98CC08803282189C8440D40CD404624",
            INIT_RAM_15 => X"9CD4E55E6CB00410842B02A7FD105706DF9E2A1FA025005632A0CC080400D280",
            INIT_RAM_16 => X"130E0174D4FB44B2C0D7A907702A748D0BA50F8FA5437ACD3B343C35039F44D1",
            INIT_RAM_17 => X"8AB3B7FDEE7B9CC735FCCE93E3AC1AAAA691AD6350E57F1F5773302B6072C63D",
            INIT_RAM_18 => X"F7F22D2FE1509BDF80E6DD7B7175B71C6531C3A86BE9F1D7A6AFD5FFB7A37A60",
            INIT_RAM_19 => X"7CA976FE488D1069D687A6F1D68A70F37CAAA367A74CBB73D3A6FFB4B1E8D4B7",
            INIT_RAM_1A => X"681A00AF8D864D8BB6D2A0916C8A9B250A76B8A977F82E8FDFBE68F8E0F8DF23",
            INIT_RAM_1B => X"BFF05FBD6AD8CA62C6CBE43BDBFD99E9EB6DD724D235FBEA9FE7D6767D811C40",
            INIT_RAM_1C => X"AF72F66DC666B39A6D66FD958ED9BC6D758D5EC24DFEBA64871D6B86D37DF1DF",
            INIT_RAM_1D => X"FBB9EB400590D7F939FF5A70A29817DC2CC29B679B2D7146BD21D47EF06F7D5E",
            INIT_RAM_1E => X"B4B15EB89456517DFF58F68BDADB95B5F764CBE7E7C7E7DF0CADB8FFD8F9A72B",
            INIT_RAM_1F => X"7BBD7F79FFE0AB8FC33758D1C1145DDD6311CF69FFFDF62EDD236FC6A0358FA2",
            INIT_RAM_20 => X"26FAFE3BE30DFAF7B9E7A5FFE4797314DAA1C1529CDBFFE9D94EB11A9F68D4DF",
            INIT_RAM_21 => X"A1FF3BE5E159FFDDEB2FBECAEB87BBCC5FCF6E23D77E4DD4C9DEBC93C10F6363",
            INIT_RAM_22 => X"2175C7B89C48CCC916D46F9315DFDECBE43E5F03D7D27F97E09E4700AA694552",
            INIT_RAM_23 => X"768008002000002624793100811F43BC315A6004052671392B47FEB7F5DC90E6",
            INIT_RAM_24 => X"8ED67F67AA66B0674CD240410F613700B8DFE7F8837F88FF4520002E4BFD7FA2",
            INIT_RAM_25 => X"7941B61372AC884EE60A372057B59CF990A6020B875C06E7C53BDF9A91F8F058",
            INIT_RAM_26 => X"8CA3CE9F24BEFA9E2BB9D89B423C327C8E050114401A62FDCD2054E166C0005F",
            INIT_RAM_27 => X"420539B476E305B8200E47DFAAE8D5D1D0724DCC3FD72C4F8DE54622A1DD1BA7",
            INIT_RAM_28 => X"EF3142B9927BEAF99BCFB066319F5BDF2EFFB11686607A73BE9CB85CF6EC52D0",
            INIT_RAM_29 => X"E3BE607B3FAC5DD39FB436C5BB7926D7FFF03EF787FF563C3FEF787919A8383D",
            INIT_RAM_2A => X"EB9963425C951C00298F26A884C3AEF0DBF539D04E867EB6FB957E817C230DFE",
            INIT_RAM_2B => X"3DDBF48E39F1AE9FC0A7CAC2B4515882877D84D415C7A00D91E87F57E95B60EF",
            INIT_RAM_2C => X"86E8AEC1EE37F6F5FFD77F204F5EBFDA614C41C1F85C32FFB05F2881BF7EB1D7",
            INIT_RAM_2D => X"60BE688D11B16D7936F4B55E0E301BAD6A96802B5719271D55D5E93FEE5335EF",
            INIT_RAM_2E => X"04FF86DDFE9FCBD3DC2A4967F492CDD5A8FFBD98573036C583F9D6D6A6138C03",
            INIT_RAM_2F => X"CE21FFE0D222852612C7A87E8DFE961BD8CF052D4757559DF3ED2417472384AF",
            INIT_RAM_30 => X"35995E3ADF9E07EB861E3035B1EF3EF935DAFFFA1F94FDCA5B833F14101BE318",
            INIT_RAM_31 => X"896B7EB5FD69B679669CBA00AA9A431956A3CE676A9D7B50D84F3FFFFFC4AAF7",
            INIT_RAM_32 => X"AA8AAA32A2C38012BFEB492278CD27651FD91BDE452EEF053E0D2912A0D49D9A",
            INIT_RAM_33 => X"C165510222E12BABC9B940EB70182EDBEEF007365AA980A2002829A05282A2AA",
            INIT_RAM_34 => X"F70811E17D8C73F1D9BEF7F7E82EFAE6C2D2DB2126004D81CA67DACC344F6458",
            INIT_RAM_35 => X"776B42A5FE80BB5AAA2A550A58904A1C6DC992952AB4532C6CB2F975BC101356",
            INIT_RAM_36 => X"4B7AE34419240F3C0170E001D6CE75F0475D5A8A9012B9BD97153AB038EF6187",
            INIT_RAM_37 => X"812017671773A9EE08641F818054455F0BABE232D2AA00081423C0BCCE1E642C",
            INIT_RAM_38 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0020203478F160F42F9A061FE44",
            INIT_RAM_39 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_3A => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_3B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_3D => X"522828280000524A124A4A7E4A527E4A106010607C38003C025408FE24000000",
            INIT_RAM_3E => X"800400207E4A0818204040024A1262124210084014407E08520A4A42424A1256",
            INIT_RAM_3F => X"A504087E764CA02840304044540424244404044024804008A40A54484448544A"
        )
        port map (
            DO => prom_inst_3_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_4: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"111F830F9851184101370588A06D3BF9AE621E7FCE632A6799C8FEFAAEFE769D",
            INIT_RAM_01 => X"EC2A08157331C6CC0E30884244916A0DE26D4D22454091290404A492016887E2",
            INIT_RAM_02 => X"96968460CA3388A03ECB45F2C4B70F1829221000FFFC7FEC346F079F13079798",
            INIT_RAM_03 => X"2251A60725008AAA056591C4000BB48C0BC29B8034A03400027B84769B520D91",
            INIT_RAM_04 => X"C13E7C640F364509212AE9CC14296E30DEA3057B35C641762CD00D40DABC2747",
            INIT_RAM_05 => X"861F8BC1993560946D92D1C0C7F046A245B5849CB751FF15B97FCD50BC7B8524",
            INIT_RAM_06 => X"E90C8E38C8E0478AD8B388F94891C9673A50BC32478E083074657E8E0EA53BEE",
            INIT_RAM_07 => X"17A24D2C636ED2478B5AE1C99D40761B1E7AA6A89DDD1BBD8DBD223E70531BCD",
            INIT_RAM_08 => X"470542C2E3C783A4C24767084C52DC209D60E95DBC096D9A0171A12D5AB99BAB",
            INIT_RAM_09 => X"5686C6CA41B2224C88D8456C1DBF20DC20A6649774CB11B69933246E9739C998",
            INIT_RAM_0A => X"3488480610A91A851E84FF08783F81AEA52D2FDC2200BC2FE81C0357FBEC1D87",
            INIT_RAM_0B => X"1620D1A60A901095D12A0973B95E20838001330138951361967847D42901910A",
            INIT_RAM_0C => X"8A370D60A0AA3E7288F4B0869FA5E703D1AE17C0EC276B2AFB747B550A8B4102",
            INIT_RAM_0D => X"95D23A0E191EBC2134B833D53D37E42B05018289A10300A188E315CE98640F54",
            INIT_RAM_0E => X"DCB42E8E77212A58842051A078007109A0D820166B8810426002844031430482",
            INIT_RAM_0F => X"C82B30679933680037A65978674DDEC2D30EEEDA78F5F2A1DEE660FFEA11B175",
            INIT_RAM_10 => X"C194E3598360AFB031A1690F4625BB628363B4C90A400E3A04DAA70DA0CC3776",
            INIT_RAM_11 => X"9DD952B29003D7767BA581A68BC41C2B16AD6EB57F1D048CD4E464190D25ADF2",
            INIT_RAM_12 => X"3B9AF0147BDB7730B4E11D9D11C1D0C3C6E0B6F242719988ACDDB17B4D81882E",
            INIT_RAM_13 => X"C653A0510A1B00C36AC88058CAC126E14E198DFB07E81C3EC1510BB08F8F851C",
            INIT_RAM_14 => X"1310B00A49902C0104004C654E0582040001103654011012021912281216B000",
            INIT_RAM_15 => X"A2E5A64B241400267194CD524499BC01D31058CD18684A817A5800B65143281C",
            INIT_RAM_16 => X"A0CC44CC94E2649242CE08191634113154562B149100204551178DE805D98EC8",
            INIT_RAM_17 => X"1AA1C248D293110CB951445117D9B6AA500F65068B8CC508BD00184F8501B010",
            INIT_RAM_18 => X"89B6054CC727D292805705A932685B6A31111371390B240EC3CC85D331813EB1",
            INIT_RAM_19 => X"316412C4900F646A36630261DA093053D98F19D2C5B653195D4A71AA5682B29B",
            INIT_RAM_1A => X"08980020680249882691A6C0488292310B4313CE87FFCD5329A64B708CAC8533",
            INIT_RAM_1B => X"2730A263DBCCAAA88712242B3BE49AA5338990229B391158C726BC7EB4ECC323",
            INIT_RAM_1C => X"F10410AC463BF80C9074917E0674A12830EFA280EBD3131E484A255D0191C685",
            INIT_RAM_1D => X"3DA2C64840C2CCE811522B42008095E5A456C98F4B25EAEA410610545024640C",
            INIT_RAM_1E => X"7888672DC999B7046A61E60810A7434450E3D33E330F321A18E8A120D1EDC862",
            INIT_RAM_1F => X"35861A00A6112A1481AF1A50A6004A05291627227FF08229B87389E08119A28A",
            INIT_RAM_20 => X"4B710C9DC948F06010DF01D880C4444BE8854062D10DD93F30A62AA7FD227C4C",
            INIT_RAM_21 => X"5BFE5CE861A20F71E8032916A78F29CC546518461522E4E14998DD54BC0E40B6",
            INIT_RAM_22 => X"40B6C18000680080125C75401AEC44E8C01A8D40D1412B25A09F7600B0C6FEC6",
            INIT_RAM_23 => X"7000000030082004A17800828F090A0C318CE120012172286317922341A2A128",
            INIT_RAM_24 => X"093E11673256B3169C12284980E92A034141E0782507800F8100009C403C0786",
            INIT_RAM_25 => X"8249144AB52CED94200A0202A88510084D938A30A34512C0CE098F08A98900F2",
            INIT_RAM_26 => X"AB6AA38578BD55CEC9AA28082C285B8C0201104838AD502AC160C13C70620B81",
            INIT_RAM_27 => X"1228D91C352915424000000AA0088F63153A8AD81B945C8789F01C86548D12CE",
            INIT_RAM_28 => X"9A22242CB58413089465B246231330D806105010035100B08761A08506094160",
            INIT_RAM_29 => X"00CC60799124A8520C08050122171281808058018C38A645D07931896B39ED25",
            INIT_RAM_2A => X"3C251301FB2CA45562245308885131119115C652B2493252340201101942D260",
            INIT_RAM_2B => X"2A086B442661015380041594608092D9CB919250100A37DDA3919A1427F66096",
            INIT_RAM_2C => X"02288A804612A2A0A102A418CBDFBA554499541660F812464011010126314289",
            INIT_RAM_2D => X"6059E332C311521E6522901852D484B423A98816C9B26A08C92368E9F8055245",
            INIT_RAM_2E => X"35188757AC5A42DEB501FE010586249AC1EA60D08F4267D2843763CFC9190C05",
            INIT_RAM_2F => X"E2975A2686A7AE0288F140141B698E2A82A835F478453A1D722CFCED12859FD7",
            INIT_RAM_30 => X"8DC6A06905054C8C36E4199E74638E6532965218A965909BA456000451343351",
            INIT_RAM_31 => X"7BB16DDB96B7845371C30B55DB96C8F6EB4B453242FF6A4DF84A76B5AEDC88A6",
            INIT_RAM_32 => X"FF7FFF7D5712524D4A30723514B2B3064A84B4742D484152FB611117AA9D9B7E",
            INIT_RAM_33 => X"0E78522BA2812C1454A502ED1A59CBD76A034756F5765DF7555F57575F7F57FF",
            INIT_RAM_34 => X"F88D5002628FFD13203066C850F10649F21319109208387641120B362124803F",
            INIT_RAM_35 => X"52979565817114DE46462844A57F7958873FC4B255C8AE549BDD1A87415D5018",
            INIT_RAM_36 => X"453FDC2219C225E421B320085A8FBFD0C42135B16448DFC226E09B3438A740C3",
            INIT_RAM_37 => X"5861917919344A4685CC0990862A11324792E761B6D41C0FCC0838C1C27211A2",
            INIT_RAM_38 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD010D2195982823226DED0ADFCB8",
            INIT_RAM_39 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_3A => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_3B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_3D => X"024428106448524A624A4A24425242522060108010543C00044A105424005E00",
            INIT_RAM_3E => X"807E7E10005270182040407E4A1252124208084008404208420A4A42424A125A",
            INIT_RAM_3F => X"A50276000854A0103840403E540424244404783E18807A08A47C54484448544A"
        )
        port map (
            DO => prom_inst_4_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_5: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"0220000000000000080040004023AD496997BBFF877B886EEF16FCF229FA091B",
            INIT_RAM_01 => X"00000000000000000008400000000000000000000000000030600000100007E0",
            INIT_RAM_02 => X"9CDCADCF90E7BD88125BCE706BF6D04AABFC1C001163DC6EFF7FD32303030300",
            INIT_RAM_03 => X"E7622EC485808C841D64B737041FF68813B149A41531A0A612FB14AE2E5B49D4",
            INIT_RAM_04 => X"C52A6A379A382C6D2F5278DA01396D0800C0046405C06F466DD18C4DD7655CD4",
            INIT_RAM_05 => X"AFE59E91BF11498940A0944996D47EE8D7E3A4EAE611AE19A965D01BA86B55E9",
            INIT_RAM_06 => X"042216E0216C85B8912250B7157D5955ADC06CB685BBF071B47D5193363C1CEC",
            INIT_RAM_07 => X"B5D49EA9D7036A45AA9E870B8E8016720C7C3102AE925262492084584942D209",
            INIT_RAM_08 => X"F665955B4E2C63DAC0078652D10120900298F7EE380092442AFD400BEC43C003",
            INIT_RAM_09 => X"D18FCFFFF3FFE7F9FFFFFFF82C0B4221214711E08904524A069491774E663F48",
            INIT_RAM_0A => X"B111114514CB11840E04828849C621392041163C00808D67223422F00110201D",
            INIT_RAM_0B => X"67459F1A8C3240FE4E6A8D028C0C088FCF471D400A19B38211004DD122212288",
            INIT_RAM_0C => X"FE2AC2A884A8CC7FBB821C851CC92B12E15593C0C020FFEE066558590E882D5B",
            INIT_RAM_0D => X"00300A8D128FA20030ACCBAFA237B7024504D36A4BA26081137F059E78991154",
            INIT_RAM_0E => X"09312DACE620656EAF24D57C08FFB14D289613DC32083803B84DC6415FD5EDC0",
            INIT_RAM_0F => X"02E84F961E3C800AC610D276182020227809001A50DDDBA3487BB6AE802BA065",
            INIT_RAM_10 => X"4915C84D6C24BAF53929814CA8A4697E8F4201145AE7415DC122A5F010433107",
            INIT_RAM_11 => X"46AAF6CFDC0791AA97B741995A3B3981E06D1A44D3711955197BB9910FCA2074",
            INIT_RAM_12 => X"3B9254954344968BAC84141C90A9C0E016CB24EDBB4D267E11775FEDD6A2FEB3",
            INIT_RAM_13 => X"0FF81FFF7FFBFFDFFFBFFFE1FF0086F3141AAB6005810A05A1595A893F9D8598",
            INIT_RAM_14 => X"FBFFEFF03FFE0FFFBFAFE0FF80787FFF7FFF83F7F87003FFBFFFFBFFFBFF0FFC",
            INIT_RAM_15 => X"5519198C859000004012AFF4FB060307C92BB732203BFDFEFFFFFFDFFF87FCFF",
            INIT_RAM_16 => X"F40B800FBA159B6DBB296562CB6220EFBE99D2776A202044D9101006FD221D30",
            INIT_RAM_17 => X"1A2955372D510AC266A5445146E27000020C320FAE1557E37154040A10200DC6",
            INIT_RAM_18 => X"111821321BA426A4FE4956B43591D1AC271E83E060341AE5F2023F0808177383",
            INIT_RAM_19 => X"CB9A360865678449975A8AE72B5C0F7BA800C1B5DC55D7D1FE2EF4EED85D00AB",
            INIT_RAM_1A => X"2508062020A0249090009252040249108806A328F4006D2AA514B42FB006ECCC",
            INIT_RAM_1B => X"17A1841358335450D4B26CD2A21B3D8F2211080B81EC040D7FA0B51CD4800811",
            INIT_RAM_1C => X"5B5C1D9D4193E40B9F492B0E0664E13AE35BE6B67AC8057BDACC155F14E906A0",
            INIT_RAM_1D => X"F25E16C87C5D0308EEC52C011514BBC13AFA1028924D0C7CE738105BD47A10AA",
            INIT_RAM_1E => X"1E1EDBBC716D44D2912B80041C44558060CFCC15955C0D600DD5E71393920844",
            INIT_RAM_1F => X"E10F8B8C100323720BEBBDEBB81DF13FF97B252E2CB4F27BA091FBD0002D1A61",
            INIT_RAM_20 => X"DB46809D15D185F8809229B150D05C8081174CA6173B99703DA466629005C604",
            INIT_RAM_21 => X"4EA47F9A7E46083716911B0D585CE937B530218E8D2AD3777EE7D3B4BC56C29A",
            INIT_RAM_22 => X"9434CCA34CC9A1CB1FAACC56168071EAC113F5265D5F6A45A098D604A820508C",
            INIT_RAM_23 => X"538D134115D860ADA57B5B868E54393B1E31E762062577697D57E8464340420E",
            INIT_RAM_24 => X"01859565800698515E10A8189EE9B323E35CE7388D73C6E7A50D0DE6739C73AC",
            INIT_RAM_25 => X"BED23D9A99FF9B77183697955D76BF0CC008822742DA45B88389193DAF094245",
            INIT_RAM_26 => X"00A85E3C5AAE2C49DDC2F6C7B013DACB319A769818A1081A7389F711D76A09BC",
            INIT_RAM_27 => X"A9C9CE3AECF7BE27C000000A8ABA95251B309A60B9DDC19EC3E391458CBB53CA",
            INIT_RAM_28 => X"32EE4CCCECC64F7E6225FC99EC64C3B6DD7DED0FD7CCEA3BF09A006ECDD1009E",
            INIT_RAM_29 => X"D6B97C86DF7D9BEDFB99E36B6658F16C6DEFBDD5DF728D6209C852C37FE67CFF",
            INIT_RAM_2A => X"8662C97BC2E8D3FFDB26D23E87BFD97E635A6560CFD93F8EED26E30C70DE8633",
            INIT_RAM_2B => X"F5569FDE08906765428FB9E6F89FBF0DEAA6064637BCA63FD02E273E5557F054",
            INIT_RAM_2C => X"4EF9AD87727C49CFE7C5DE942B72AC7F6D97DE18920777FDDEE9EB11122A4E18",
            INIT_RAM_2D => X"A1BCE33AD2D8BE40A4E5BB7D7BBEC2CEADBBC8B6F87A4A56FBE0B891DC57E4C6",
            INIT_RAM_2E => X"E0948817C496E9DE8EA1F88F627B7460106691CC4526DCBCCF2CD2F003733C4E",
            INIT_RAM_2F => X"0C840083AD485153ACD3C035591630199B8C096CE4DC557D6D55FCCD738573D6",
            INIT_RAM_30 => X"924C10EFAF3CB9B62486512344C61ADE6F15AB67F335A52513FC85AFAEEE8400",
            INIT_RAM_31 => X"EA4C912568003BB493CE04FF086C188980052BF6ABAAA2FD5D658000011277EB",
            INIT_RAM_32 => X"FFDFFFD75F145247F03A0AE7F1E1EB2D5A99D2444108C6A5CFFD7DEA6ABCC241",
            INIT_RAM_33 => X"02C12B12378356DE2C52041CA7A320C51E0D7CA9F5D575775D57FD75DDFDF75F",
            INIT_RAM_34 => X"6CAFF2622B8D518F63C6030424188FD357718970D25A30CD0731E532DB23002D",
            INIT_RAM_35 => X"D2F8735647315839EF6F683C64773FC73464D5FE354936D50823A5DAEBEBDBCC",
            INIT_RAM_36 => X"59BCEFFBB68A6FF529B3B0D92970010BBB6C7D872421210E190E1CCC47A485EA",
            INIT_RAM_37 => X"5B438D714D4E3DD115E8BD1286EAB5FA1D71BD8F4508BD4BDC8838F9D27B5522",
            INIT_RAM_38 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD894D29B9D3ACCBA3F27D9DC9911",
            INIT_RAM_39 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_3A => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_3B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_3D => X"020028008000524A024A4A284252446240001000101042000054265C7E060000",
            INIT_RAM_3E => X"8004420800620824402040024A1242124204044008404208420A4A42424A1242",
            INIT_RAM_3F => X"990442000864A0284030400454782424440404007E404808A4005448387E547C"
        )
        port map (
            DO => prom_inst_5_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_6: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"FDDFFFFFFFFFFFFFF7FFBFFFBFDC0A6DBE6F8CFFBB7FE7A39B3DFBF3BEFBB679",
            INIT_RAM_01 => X"FFFFFFFFFFFFFFFFFFF7BFFFFFFFFFFFFFFFFFFFFFFFFFFFCF9FFFFFEFFFF81F",
            INIT_RAM_02 => X"B607E624499300E4DF6D95CB62F62FB75403E400EFBC3BD34080FC9CDCFCFCFF",
            INIT_RAM_03 => X"C9F7627EB100872A52FB5141D65111E6C8DA0ADB6CEC6005C61D0E366B20DCCD",
            INIT_RAM_04 => X"4C3838641E940623ADF28CCA14BCC07104C112BCC9032C48E925594CB886A604",
            INIT_RAM_05 => X"B657485DCD62AC0662C8C005DDE7494C9CA13AAE3234BB0EE1B708A23A2F48AC",
            INIT_RAM_06 => X"96632C3232C3974CDC1172E1779D8C6738251819975DB8146067301E0C0277B6",
            INIT_RAM_07 => X"0776C62C316FF94B0BC3A0288DE6A62B14D6C1A2DADF9BDF85B2CCB02CE1DB2D",
            INIT_RAM_08 => X"07B78D38001FE67E56CCE399DE36D7DDBD699D5CFC5B6D7A1421CE06FE40DB6E",
            INIT_RAM_09 => X"9693E3EFF8FBF1FCEEFBCF7CF9BA6C37640DDF7FFE6187B19ACF089D4C038F66",
            INIT_RAM_0A => X"7CBBCB2CB384BD0D92ED105D0617856E80441124B31DE58B8C001607FEE66889",
            INIT_RAM_0B => X"3D3CF1BE8C84DDB000565880A776E5C0E13166E49F47119A4CA1311CF97B965E",
            INIT_RAM_0C => X"7EE296E8986E64C6DCDDE59436641567648CB84DEB7D7937F974F038D838274F",
            INIT_RAM_0D => X"1889D25CB816ACC6627802052C61A4099B7B0EC923971DB3B9F9204BDBCCFA45",
            INIT_RAM_0E => X"7D361CDE72B925658DBE1F7C4707E195C5C665B8118C3C31B196C261DA85A5E1",
            INIT_RAM_0F => X"1C5CF062CA6F13854A59BDEEEA07E3C6559EBB3618111895CBBACCBCD512B5F0",
            INIT_RAM_10 => X"2EB0B348C0B62337739B1BC73192392592C84E37B7AC141CFE65EE76D83CB083",
            INIT_RAM_11 => X"1D77401A0C0CCF5DEEE561F7F7E68CBE72E48E570B047C772CBACC33753080E3",
            INIT_RAM_12 => X"19B9466E6D7B527565924244B20C5DA22B60D21B6030D9960699E11209699604",
            INIT_RAM_13 => X"F7F7FDDFFEDFF6FF7FFEEFFEFEFC4E51EC0888848E1F2046347B66608D8A3B39",
            INIT_RAM_14 => X"FFDFFF6FFFBDFFDFFF57FF7F7FB7FBBDFBDFFDBFF78FFDBFFEDDFFFDFFFEFF6F",
            INIT_RAM_15 => X"CEEC06DAECB0001569589D5F267AFE086C8FED5DE41DFEFF027DFDFF7FFBFBFD",
            INIT_RAM_16 => X"BA42813453FF4EDB60C6BF8DB6E267BC56CB69BBCE636CCCB3B2B4B103CC46D5",
            INIT_RAM_17 => X"881331ED7AC4EFD38DFACDBB236790005719AEA2FAECCF0D126A30A27562C61B",
            INIT_RAM_18 => X"CE618EEDCFB393738178C476C36CB61F71307F6803F677575763DB2D8C3118E4",
            INIT_RAM_19 => X"36DB5B7BD2850018CF936621C6863095A73F7BE7442CB13310B9C0BBB96EEF16",
            INIT_RAM_1A => X"0408002024010408824080002008091482ED5615E40012EE630C3B2CDB2C13A7",
            INIT_RAM_1B => X"4A3E508B49DC6BEAAB4F3F0CCCF6D8F568F2DA00EB384A7F5324932319800010",
            INIT_RAM_1C => X"2E43664448EFF19872648DBACEEDB76E26439BCCEF2DFBF664594B04FBAE72A8",
            INIT_RAM_1D => X"3DA139003D7A86B2F878DD99DAFB70DE1A19F3FB7DB3B8EF2633007664CB1999",
            INIT_RAM_1E => X"EFF4FDE394D0E19B6FD89186C23CF071E6F1CC8F7FC4F1E48756B0DCD8ED6D0C",
            INIT_RAM_1F => X"3C766E63DB6481CB39BC8C68831C724633186CC1BAE9D608A5DEF0FF219C28C1",
            INIT_RAM_20 => X"24C921BB3332DC66D9C1706B6C5903129639A3BA4088EDB496EDBBBFC2CC40B6",
            INIT_RAM_21 => X"FF7CCCEFE1996DE3ED6D8CFBF1871BD98EE7646242664EB2E338BD0098386371",
            INIT_RAM_22 => X"63FC93ED92CA4DC61B01639318985C88F01680E307C42311C0124700B28BF9B4",
            INIT_RAM_23 => X"414D536A41D144B6C4624A2B00366D8CF6734A4A2DC465B308462CCBD1BF9CB8",
            INIT_RAM_24 => X"CB76E03779E019E2C4E4028219C38C202C9384E0D24E569C2E4D4D60B670CE37",
            INIT_RAM_25 => X"E1265727652C8F0C422BA8C28A0FBB893B0881E00403DDD8843B2D8EB929D0D8",
            INIT_RAM_26 => X"C228A2050470925E29A35D8D06242712CD25C9241898204D85A710947C802013",
            INIT_RAM_27 => X"5F9CB25A3631964C20007FF5754FC631A97D4F93986C30CF24394625658DE9A7",
            INIT_RAM_28 => X"C7E1B221EA10E38F64EF31CEBF3368E1C712BB1B33781134CFE54C2123349A6E",
            INIT_RAM_29 => X"7DCCFC5939C4EC79CF0E1CD43BA7AFC716900A21BDB9DD0FCC7ECE1063238407",
            INIT_RAM_2A => X"499D7BD86619EE5574CD27C80D39F71E653FDCF1B366737233CBB98D1E7B330F",
            INIT_RAM_2B => X"AAAD6B6AF36195DA637C6EFA3E36E8FE97FA02EC26EB46198AD8DAD8C11260AF",
            INIT_RAM_2C => X"C23B9D130CA49818913D3A2C1FBF71C5B0C774336F903C677D976189D98CA127",
            INIT_RAM_2D => X"CEC3000F432029B3FE3F211712944CA54D1940F193204C199C9F49666BC11B38",
            INIT_RAM_2E => X"2F3982C7BE09AD4A32196807648A2495ADF98FD2B15E604B52F12FBBC811C953",
            INIT_RAM_2F => X"E33CB578DEBFAFAEDFD530DE8FA1992072F31B116644B18C72F9F44116C79ADF",
            INIT_RAM_30 => X"7FB1E62675F7C2CBE01032DCA16BADC570C1CBF7ECBC4E7E6C5425D4550BE1A8",
            INIT_RAM_31 => X"59F878FCF5689FCFEF34BFD52FA2422A56A3C113409F7813007F8D6B5F80FE9D",
            INIT_RAM_32 => X"00000008800AC11D556264251ECFA68C056FBCCB040C614A0240000300D2F6FF",
            INIT_RAM_33 => X"C744FD00E1A7F9E9FBFE4777FD50ABD11F0E57FF4808802282200888A20AA880",
            INIT_RAM_34 => X"57781E91788044213E091339886F337D0612CA646CD48FC58EE77EDD7ECEC466",
            INIT_RAM_35 => X"662FF5DF9CB107BB23A39EF7B95E7372200448DBDC18F9C0DE0EF379BF494806",
            INIT_RAM_36 => X"06F6612D770080980A40D293FEC069F16CB2164CA033C539F69B37741AEF1CE3",
            INIT_RAM_37 => X"0100046606572583002086010800054C0F2DE8371AC0000A9003E024840C7C08",
            INIT_RAM_38 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000C02060C000C0DF50F68A580",
            INIT_RAM_39 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_3A => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_3B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_3D => X"0400000000000C34023C2E302464003C00000000000000000020460024000000",
            INIT_RAM_3E => X"80084204004204423E1E3E02247E3C7E3C7E7E7E7E30007E3C7E7E7E3C7E7C3C",
            INIT_RAM_3F => X"4200420000441C443C0C3C00480018FC387C7C000000007E1800383000002048"
        )
        port map (
            DO => prom_inst_6_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_7: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"92225124929249248894408541300A6DB00792FFB12FEF240371F9F190FB007B",
            INIT_RAM_01 => X"0422500891088848884109240412044442091020842411042041088241144552",
            INIT_RAM_02 => X"9001624489A10045D16C944B02763FF55405E400BADFE5BFFFFFF00000000011",
            INIT_RAM_03 => X"49F30426B100842A12B25160D6D991E6C8C81AFB4C64400542140A342020D84C",
            INIT_RAM_04 => X"883838649E1442A3A1F70CA9094A5AD4A52D56C5D80CAC58D9645944A2300915",
            INIT_RAM_05 => X"A276585D5273AC87206840415DA74B4E9D213CAE3234B308E19608AA38250844",
            INIT_RAM_06 => X"B6E370363701B41848117683379C8422102D001BB41FB8248067301E1002C636",
            INIT_RAM_07 => X"84724A241226DB4809C9A1100DE6A63984D651A2624A09420496DDC12CC10964",
            INIT_RAM_08 => X"4C3C8D784218667F524CE209881213DC91099C14744901620044C802DA414966",
            INIT_RAM_09 => X"169808000200040100000002F8986E37654DDFF88E20860382DC089D4C239F6E",
            INIT_RAM_0A => X"1A55A50C3384B549B64C381920140D4008004020B119D4834C10064000006001",
            INIT_RAM_0B => X"0D1C3E528444D9B00E561C40973AE1806031C464834F03D34A11233A34B34A1D",
            INIT_RAM_0C => X"81E08228382D54C298DFC59535528176240438C9AA757917F95C7428981A2647",
            INIT_RAM_0D => X"184B56183004204267600220A061A004893E1D609106BDBB553920A011AA5AE5",
            INIT_RAM_0E => X"2DA65C2472B824F109BC594C2401209C01A0E59830002C73B396C6015B85A163",
            INIT_RAM_0F => X"101CC0024A6C32005CCB31908842211604D8B326101118B54B188CB4D502F5F0",
            INIT_RAM_10 => X"0BB04344008422327B1393C43396A931B8C8C87227A6141C0E2DCC76D830A082",
            INIT_RAM_11 => X"102B400E8004C40AD6E4614466308ABC7165AA57060A3A736A188ABB300200A1",
            INIT_RAM_12 => X"19B4C2CE666052C0619246C4B2245DE02B4009000402001E1051410804201E92",
            INIT_RAM_13 => X"000010004002001000200008000AEE708008880C86112252345B36C0048833B3",
            INIT_RAM_14 => X"0200080020000800200008000800400040002004000040002000020002000801",
            INIT_RAM_15 => X"CC0E00DAEC3000194A52B80C606262092D84A110241000000140001000200080",
            INIT_RAM_16 => X"10438134E31C28000400B18422CA60FC42C9C03F066366ECBBB010B00B004807",
            INIT_RAM_17 => X"881B30810845E6D18622EC9B6236A000030986A4F0644601226000A2F020C403",
            INIT_RAM_18 => X"C4C088B1A9B24BEB0178C4D6C18C3C5F72B07A28063647CC4721026D8C711864",
            INIT_RAM_19 => X"07D901787004001C459326210CCE00C6AF707B84440C313B10B8C4D13B2C6E06",
            INIT_RAM_1A => X"00800020249004081008924124080914000000020BFFFFEC638C31207B6C3214",
            INIT_RAM_1B => X"CB3E518948104042F84F1840401018406877D800A00000F5122597005DA44110",
            INIT_RAM_1C => X"6E436E644CF6C8D86F124DA26CE9B66E2F46BB466E2CE068661B4B05F02F7D00",
            INIT_RAM_1D => X"202139803D3000B2E0209DB9101160989A5916381001B0446631006064DB1B99",
            INIT_RAM_1E => X"C71478E35468600B01A93082C63DD073AE4181844449C08D8D56B0DCC881251C",
            INIT_RAM_1F => X"7C762E21DB2481CB6BB88C68811C76C63B18ECC1BACDC6110DCC70BC20940800",
            INIT_RAM_20 => X"66CB633B3376DC625DA8A0856C490392B779E1BA4088EDB4A6CDB9BD46DCC0B2",
            INIT_RAM_21 => X"FF7DCCEF40196C8381658D8840043B119B86A46247665810E2203000141023C3",
            INIT_RAM_22 => X"3124862592C0CD0F07A27A111CB80A48808C7C21C205029100010400228BB3BD",
            INIT_RAM_23 => X"C14D536A45D144B244C24A290076E58CC2E64E4A2DC4C5939C4C2DDBD1B918B2",
            INIT_RAM_24 => X"4B72C08871D2413188E4829219C38C2025920480D64856902E4D4D60B640C833",
            INIT_RAM_25 => X"2166D72DC524870C422BBFFD4808A7016B088DE3000B853800336C8E9968C19A",
            INIT_RAM_26 => X"C629E6050C619658692170C1022C2232C965C92C189020C70587308485891032",
            INIT_RAM_27 => X"1B9CE2DA363196DC20007FF5554FC631286DC716B048384C26510685218DF9E6",
            INIT_RAM_28 => X"03C11245EE31E38E6DEF2188BE2068F3C716E10317783020D8EF5C256774BA0E",
            INIT_RAM_29 => X"7D8CDC0131C444798F040DC0116E2C4336B0166109A15D1FCC7EDE31EB238622",
            INIT_RAM_2A => X"4B987A78AE1BF80005EF370C0739371E0D3E5CF1E3677332370BB98D1831B30F",
            INIT_RAM_2B => X"0001022EC10015E263787F7E581EF83F062200C626EC4E19021840D9C112400C",
            INIT_RAM_2C => X"C23A8D170CED981891256A2C1D9B31C0F040202103900E6765976089DB8DE16E",
            INIT_RAM_2D => X"CFC3000F43632B49C39723270C604B184D1940F1B2A04459BEB088666943BB38",
            INIT_RAM_2E => X"AE6302C4BE6BA8C22A084803225A0855ABBBC528B1DD122B524A8D33C1209153",
            INIT_RAM_2F => X"873CB568FC3F09080F4400DAC600092017210911A6081DCC4979244124815884",
            INIT_RAM_30 => X"7FBBEC46E8B3CAEBE0100275A1092081D0C1E5716DF09CFEEC022D800529E1A8",
            INIT_RAM_31 => X"596CD8B4B568A4DFEF3DBF8027A3422A56A2C003E514582104BF8D6B5D80BB39",
            INIT_RAM_32 => X"0000000288964258156302504F5F660C054DEDCA20CC201A0206160601E376C9",
            INIT_RAM_33 => X"C7C57F084106FB3B8B1E47463C0088D11104F23C180222A0AA22A22882A202A0",
            INIT_RAM_34 => X"5775469089F04C623E19317B486F653C1C22CA642CD685C10EE47EDD66C8C226",
            INIT_RAM_35 => X"763C75FA1DB107B865E5B8F7B95E77F222244C6BDC1879C0562EF779BE000946",
            INIT_RAM_36 => X"06E5AD6C882882990A40D293FED064710CB226CDA0330D7B189B344442EC35E3",
            INIT_RAM_37 => X"03020CCE064769B15020A6030880234C64E9BEF8E98A81489083A026140D6489",
            INIT_RAM_38 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE8840C02862C088C36E19CF1D315",
            INIT_RAM_39 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_3A => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_3B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3E => X"8000000000000200000000020000000000000000000000000000000000000000",
            INIT_RAM_3F => X"3C00000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => prom_inst_7_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

end Behavioral; --Gowin_pROM
